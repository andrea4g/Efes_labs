��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F��J>�����>�����HU�k;�� �[�+?�w)݁)��>7Ý�4�B#�"u�%��R9�*2�	φ�v&�f�UxJ�%�����OOL�mF4O0��%�O6?][��W5Ff�i�]�E҅u#��Vg�n�����g9�#���>rh�W&��zCu�M��{����,l6�`I��3����
X�	�@�#��꘲t�}p�ũ�g���.�pæ�dbB�:�`�(8����Q���E�m5���[\[��Z�Xe���z��e�ّ̀�4��'͐??�r���4U��e|{��s�_
���^��5���ЉS�u^R��r	
 K�Ԓ#tO���?�M�ΟuD�(}�G���|E�,n���;��"�z���+�rW�t�ǟ��[�z���Q��Ƈ�b]e}s�;�H�:��(�=����ݺ�����)%����j�⽾I���G6
�<=h��/�[m�S�\I�.4�A�1��S�S��h$��Mj�1�~�P|ul�P�,hM����R2��U�&tˀ.?���9i|������u��F_8�����-�'zx8�~�$	�	+��D\ߍ�b�+/n�f i��O>U�9���mx�������V�K�`?2_�ĥ�3?@A�ʺ*��P �j�C�
����ï��b�A����[���GE��\
���k:
�@�fv6�xR��G��� +�U�.?�T�:y4�_,��7�&��!J�+9?[X��b�1�#���l��;�l���@�7��-�c�)��(�E��V|��i�P/��0��9���E��bQgb
�fYR�E���Do5�����6�r��"�Ҝ��9�=�N���5�Wؒ4��P�bЊ&x�`
'�97^�(9�!W���Dxp@p-/��0Iﴓ8�Y���v-qk��;�Ң7ժ��ٲ?������TH�A���o~��pI��<C�@}|ل1�ў%hz�&��-p�n5�,I�)3�����*�}{�.�O� qI�naG���"0Bσƥ�pl?[� ���,.χcFP��&�?uP��
����������K�,��hXJ��Q��^�M����ϕ��< ������h+ycmh���I�s3]��6�  9UĿq�����⨼�LKU����,��#(w����[L�ޛ���N`c�c x�j�Z6l�iq�ﴌ�P�	�:M����#Mt	��(4Tq�4p8%�;� �o�;*�;OI����˲n��>Yb��EL||;�Yź�>-VRx^$�S���/�]��{n�BX�'i����f��#��:^�:a�:����1�./���)6sm{z�e�r��?f8�XP�796��ߑ�]x�jg�o�۟�­x$_����L� 㲔?��r��t`j�{Z^\�L!����k����S�{i�z��n�ӡt����&��KigS�a�_w
����Fu����oe�k�XVM*E�pbϛ=��nۼ��"Ep:�����*t��Z��k i~#.��`���A�ȋ;�u�U���'y��ʚa�8n"�f�&��Wqf/��D�4�8nBmFr��@���������
��|�QM��<����k�&�di|g�ᄌ&���S��=1�'�:��[��u�b7��jQ��ݼ�@���E��k1R|*�뚩�޶�(s�.^Z�B���"'�dk����]*���������H����H��M���LL<�[����e�
"(�h$)&�����Yz�-������Wb/�H/��<�'�Z�L���2����q�LL|�ǖ��0�q� f��!86G�l���#S��G��˳���[i�׉� =��E�]�Բ�}^�i��z_�ؤ�"���������;s�=�o�W��((�h�q%���T���-l���5
V�$���e���@�D�N�2w�Kх]�6ʌ�(� (�W{Q�x�Mf�EpeÜ_�)_3>qM��aR�ɡR�:�HDK,�#�hu��5�~�����⺰�Zz����:��Fӥ���mL�&� h^�͞�M93�mh|��C��M��o%��.FɺH���p�Lz�/����[�]���X����Ae1�/_���U�K*U7?�6� `�Y�ԟ*�k�OJ�����3L���ĺA#���P�B ���C+
䲑��;iN���A�%s�<ḙ���=2�h�o	��R@����r싕��[\A��'cq+��k�� ?���7�#շ L<5KL*�yA� �~i�\���D��Z�ǜY+�j=�%P ���gy��
GR�HU���I��gY.�Ǒ�Cs=�HW!hV]�\�J}��}O{����\2���E7t��ϟ�q�\��=L��hQc�v�
��H�U<�����/+���S���v�e�c-7���Cji�-^��%7E���7�W���N�pA���I��}���p���dY]�Ƈ�g��d����g<�
C�Ǻ��ͮ�.���;�~hK�}վˊK�A�^�ah�u��"	�O��Վ?� �5ɠlR � �lgo<� A�_U)ƕz��E3b����bn���.W��QhWK�A#�:�U>��g�
�DR��]��`�|��J���#K�� �cj���O��L��|8�����q�U-Z�#PZk�5ײ�:k���tP��x)|�®���6 �!t@m�Ao��<�A�.�s&��!e��\��x�8��i�6n�����(�Ο���V����/ֻ$�`�Ҕ���� $G&��aKD��-IHj��� }�L+�0����oi�W��vLi�͗L>L���ɸdol�q��A8j�+�Pآ����fC1N�	��/�=Vn�{�P�58쀲���$8�W�:Yl#�kX���ڿɊB_�ڮF�Uͻ�$T����z�@9���'<a	��i���)H%1D� )�6��8�Lu2u
�{�[�k���
ߘW��irM�BR!?�p#�	��Sx9��53;����h��i�饧Y������~�zA[�J`��O�:7m�Q�°\�����Bo��Ohi�d�(�A/��kw.L)�+p�K�u�Ƙ��@H�1�����N�m2�P��x�t\�.�&�puĚP�͌��R!��5�?����!4I��2��&%1���{��e��C�ԝΈ?��o�l���Xٔ�ڋ���:7#�ڸ�" W��'c�ӄ�h��'_�.z�Ϙ�1�d���T����+�q%�?�Zp�]t8������x0��N�M	:��3/�wz���L�&D��?��D01���ϙvIW�)_�F��F{���Ҥ<G���T�P������Y\�)��s�i�{=I#+M&Y���!"}Y;�J��z�܉��e���2�o^i�X2���_+7.	�^����P��3�t�r6��]|�ד���xC��0�o�̎mи��Xf��d�y�'�8񰤫��<�V)U��9@<fv�4V�QE�l�mT��=��E���UG��r�1�b� 9Z��e>����F#$�z�߰⏝^��O#��IS��cք]\ĝNH�d4۪�잼��B�Z��L6���x�M=�5�������������E��=daq�q��$x�҂�d�@��%<����	�y�vD���yqCdvu�I�>
V��6���|�m��הd詉�f���ԥe~�O��-���O �����$�L������kC�O��edy�tH���%�N�놮'z�Y�,���ᛲ�� �
�������C�^E�_�b��BK�ל�{&�Gt��KD���и���m����Ny��U��4J�l�E`p��{�'�Om��d�<��=�+�����Z��`�\&V�ͦs`ш獍UR�[��������Fv�֓��K�h�V
jK7�(D���l�.	@��p�9F/��b����uo�,V�L��\=ƛQ� �ԗ5���G.㱮�p�߇��l��jSe|����{�]Fn΍�m����|�����E���zR�')Z|��S)Y5eD$p��M$����&�.����p �[Jܠc�j�u��'~]	t���"���Ł��Fp+^�5:�b��d��:�A]D�7��C^��~mo��_|�\�̔�'�+w�թ�I������^M�J&�����/vQ*2YS��4Apk&���@�)��c׸�"]���r��q��v�o6��*�I��W?����EW�}����Q�yr�~�,�竣+�.�E'�vjC6b�x@�q��{��g�r��Mzl/��
�B�`cC����Ya�w���z7��!{�G�X���Z	�]�}bQ䔺jk�3,
���?���A�㲈.����fDC)�k�����tݠ� <��0���+g���=�
<�U��CA�m&�G[Ck���،�y�������3�#�D��<��X(YI�b:���0��A���13�Gb�ك�2-�Ng1��	���,ܥ/v-K%�"Z��6���f���հԋG-5m�g�؉�Ҭ�ڐ �td�!5�E(.᜕0h,�L$s��]iH6`�8����~�2z�^6�����Q�zXuu(|l�6zͼ�0�:'�낾��W9��\�q���g���O٠�n���|v}�商J�X�������r�,�]x4��b����J ,���B�o(B*\�/�iD΀%�]�8��_ӓ�I�k�f�!��5 �>-��������]���F�,	�1-U`��T��ۉVR��#��<e�'�g�	�8���;�~y��Ķ�iа��>��ԍ �5�p�s������T�����\O���o�[_�w�ǮȻ��q��U����(#��GP��l��`�r�#I�#?|��g"]V�"�0/$�"�K�Y.^������������[�;*YaA���޵g�Y���0�!�X��h�b���t_ѣ �>DIMz����\eM��@��]�^;��U��L�}y��[���s.���a8^��u6�'۩�ȏ���^'qz!"ݥ�G��R������"n����ZV�R�瀶���Z�z׷��0�������������Xl�wi��~VK�[#v=!�2ps����A�ʆ�=J��f7�6尺��vυ��̺�^��s:���͝p�]���E���KQqL���'ӓn���4xR������Ź�$�k^MJ�������F}TbFHX��>�|Zr��z�Xa5����z敺�Q�[��T�?&G�ltЏ�bpɺS�<p$ƭ\�g!�����鴒���5��v��
��]߲�ք�/�P$tֲP��p2 ŉ@�,� ��8�v�Am�.�%��m^k�F��́Nb�t��?�vJ�T*�̕.J5��w"��|�AËl���\��:6�kp��d�/a7߀쁰	���2��씲��QQ�#y�`1)l��!�!���x������Ȼ�kQ=�h�"*+J�d�^-�|�+!�^LL`x$�Z��4L���֊y��h���Tg�Q���οD�}M ����c+߬-`�$����J���|�i+���1�7rTG�H�C�P�!�����G<��������	��\�j������g��Ln��)Uy;�"}��1���^8���npY��2�>�Bc�����}�mt�@��.��J<럧/�5��Q����4(�֟�N4���|&��6���s=�:5���'�b�����
"dJd�K�yQ�~���bWL��s��#��4g^_[���"�H�Z8��%c�n�Du�ы̽����iq���b ^�iBqǡ��8�ӻ*�NV/Kz[�r0��?wQ�p��<�1��9S1l���j>�M�*�H�`����<��n�p�Q�I��2���	�0���8�����Dm2��,X�χ�۶Dk�2��4�)��n�|�^[��������n��u���� ���f<�8F9��rv8�:���~0�
K���C������$�\���E]���-$Ea1��&5���L�op����ʮ�����$���Ӽ�"ܾ
��.���N����X.��K�ꟌI��ޘo��K��]��x!�4͔P�;��;�c%���!�t��8����N�)��iFV�~�Hn����Ǖ�Gi&�{K5��W:!>Y�4�D���v�_�Hz�r،�f���K#Vz'OG}xm������T]I>�8S*{4�t��Ps�h]�c�ݹ����@K}P-N��A"JW������Z�pj�n�Ŕ�u�bc�IT��.X�o�c+��5;�_�h�}��.Y�y�.U�S�i��/?���Z�+���륃��C��Y@"��grE^����mI�d�O�F���oHO����3eIuh��
��w�=h�� �ƢK��,�g�
'.�JC��3(�!��̎�;�s�WZO���R08�� �o��cl79ܘ�U_����@k�E��*X��e�Ā�
ɖ�l<��i��e����äup���{�3Ec�v�J��{�X�?�!!Zŗ�d1A�R��N��lj���o�l|�
,jЁ�.lP��6����!��
�J$��"��1��^lR1��QP�g��Yw{��鍖O�����U�J�����S_RC]�"�X��s�C�9cIW���m�i�9���Gko��:f�1�dSƏ=61�1w_T�×�J����aD�H�$�BP�����w�z*�Jy��0�s�,}��o��K�3��D����<=.4��`�Ʋ���hI4��)y}7���5~���(��ם�����,�|�ȵ�#[�#NG	�,����G=�M��2��=�K0��T�UHD��Fڍ�����V��v9Y7�\c�"�4��q�"�i����ۋ�Y�9��۩{�J��P�s�94�*j��5��u�|�PUpB�m�P� +n)V&��%�ӷ�����2�`��t��c៤�+�&��v(o�G�Op$�����
r¤�o��}���d��k�7��ӿ��vT�,.�xE�0��C�8�$J��d/g�t[ �SG� ��d�!�I����W���a0��K
�T7�X�x��[&�4�$:��,ʑx@����Q�͕=lQz{���|;�B�Y����GK���#k[¡�"�*����z����;fz��H�sOXG���4�
�����l�m�A�".8Yq�BqD���� C��q��"$]Ɂ����dݷH3|&+X^��:K0d��&GG��D}�:r����%`b���z��0rgvr��܉�/R'w7��$X-�u�V�yy�J��bm~�R�'q�����.�'0�^�ԕ�Q����g�u��K\'����1�g��K�����]�=�̎H�d��k��d�����DJ0��u����hE�X�爕i�%$�8`U/��[E����f��G��~��*c�����m�7(��`����X�i�j�������N��UJ8��q&B����
#L�� q�H}{�UK|��\ |Ό���oH�,0��|�p����NQU�� �IҼ��뽇G���U�v�-��,g6Y1����W��ڃ:�"Ǻf9��%�wT�X�'���˂"H�\����H�NV;!i���u�)z0���a�ia,���N��������|�.>Գj�WjB�m]V��a<ZU���	�NQJ�����E�Ѫ����O���������/�o�}���={�A�I�ܰ��h&�c����'�wHt�p�mC��:|�Q:w38+��q;�r� Sg���1�RC�F��?f���4�d\�B��t��*{0M뷰L�n����V�$��tv9� �(<����.}�r��)X�]y^�3�a��e�@� )�k�>�#ـ���J^�X9��v�d�΄�.�ֿY���c�c�|��f/���%.2W>�D�R�[T��_����'W5�d��T�o�kC�B�_�,����N)O�T�4��'��1bz�Bd ��}~��u�i�H�r��z�I�7�p�!�JE�~�^>����&ۯ���c�{��-`F�#�x�)z����#��J���WH*[�s�"������u�vͱ�ko�P�)����FA0mŢ�6t�0���r���Gn{��$�s��@�Ta��q;�W��=��[$�ָ��@����nA�ht��!"�3m�xD�P�RՅ�9�la1%̯�(4�C�l�|h��ih�?G��(v��[��k~���=���c�. �kG�\Y�R��"�O�����g,���Cm0Yk����=����H��g5������xk�O��O�L�d����
m��]b]qi�=��U�Z>�M�����;��p���kQ�������6�-�n��	SˊۑH���=k�"OO��8X���Z]�a�k��J��2�	Ha�3?2�7/e#rk:s͠�Uq6t�1Ů�;�������꯽:00�XqAT�b�O?*�._�(�5�C�t���̜٧���r{tѤ�=`�ZVsk)n!kkk��񯩕�;��$��z��@d�pȔMVޠ�a��#���u��IC�mSS	�U���ǒM�X[Rؾ�~�����;6��8C�9�=bh��᪉�/�1��c�k��H�+��2r�w�i�4`>�FO~10Q^(�.�l�%2=�~g�i.��ߢ5�^I
E`,���	��l+���|��)����O�X��^S\�d%��%p
��0)���r���Ϻ?7�e�ő�i�s2���!칩�އ�v-x^��$G>?�>�-cAn�|�AhQo�elC�W,cC=NH��,Yg]������r����k�+�N��JbR��)� �߂U.���l��i!�C�vS�.�Q=����v3J�ȃ{&��7{�@b�����~x{'QiE�&��������t������*Qo����v2&a�E4�(��_�DM��[��ł�s�p���0\�<
�\y��K���}�<HH|V`����yg�<����e{�Kt�gV����g�k����ĵn��"p��͞藃�1(qc�51&z�e�eG9�k�Ϙ�½G�Mn��5|������O�\��tÿA�b�@�&���I�TY�$�Z��\�h�� ^��]qrH�����ȳ9-ȇgldM1eS(�!`�q�Re؊=���u�k�g�Z���>`�:ȿ�����č�p�U�@�_���+%*o� �Ͷ8�p�hBwh�X�z��P�M`Uri�ur��}j��jkx+n�돘��V;�(��r?,L��t��^ݰp���5�i#����q��8 ܡ 9�o@�d��:H�'W��d��`p�2ڕ�-����?��V?�z���R�Q�ٔ��1a}kS��u�w���i������������p,��yo�+�''� G��U
$4EPU7f��ʪ��.�Sp�a��	���`%����d>�iU����^H�}���V�Ռ�Jco1đ�8����4��|�$ߔ���	��|��v�Ճ�76Q�OҀ���ʓP2N$YE�wj�G�M��Dߙ%:4��<骋=$]o�?��k�x�SKۏ���څyQ���2�D����3h�,Zb�(�oO���!��C\�*���4��a� f��)���T}�Jg�*Ŗ��N�5�Ӭ��=�z0����=pbU�:,L���(�s�v	�hS���U�ȡ��ҹa�o�(�a�&-zhk�s(h����<sԘC(]�M	{�(�����zF:���&[{��4<H&�I�Cʿ<���C��_VN.ov@���plc�r[~��:����:oƮA4J�%�*?!�����#�&�D��T��9���uj��3\���IS/A��E���[��lSV�P)�K
Wp���Y��3FN�8&`�ק�� 4`�r�7i&L7?�Pˆ2�oȺ|�1�r':������cv�١��@ �m9&Y�C[�|�%L�	\�(�����N��G�pVnY��	����>��.�D���\t~�L,��n��;*����<?�{q����N]�?@}?N�3���x_����|��S<̝j]�s(g��|qE8��Z�4U�#���s#E�W�bo✒@落��Ĕ�j����ۡ7yU>Q�%��<LT�+z��c�ϳ��Z�E�r����P���z\�:e��0����	x�T��oɜ$�5P�i�W�k����e���q&��(.���l�8�ﯪ�khq���H" ���o��q�N��)x(.���xh�[+��Jf�A'u����`�__�z�/����ˎ4G�r�C}�|����Nt��`'b�����G�85R���v�m�� tJ)�]\Q��
`��"��y���r���h�]�w��՘�������C�3�L�w�W��d�4��_���om��n2Rr*hV�|cį�E.=�R{�{>lm�����ƾ��y43�A����
�l���+Re3�N?9�7��a�O���᫪^f
�^p������V���]�ߌ)x���@�w���d �����(����t��uGSo�P��Ά0�dO�I�;K���Y��z��]���ljB�g��A���I�(ٍ�,y��� MÌ�'�^��U�d��E�`�I��7���d�P��	B�|��f}�=Q����ɞ3���2�Ĉ	\�gy�J�;���gz�k�i+Ӯ�����u�l<U��Ҙ�Mx�*��~շU}�mJ٩Z���=<]�~�/���_j�jW�7�v�����I��Se����Am�](C	0 �ik��'eA�_���{�p���?o��\��0���#���������j�=�Ė������=�""M��Ҋ��E�j�Z��� ��$0�D�Gk�(ʘ��j�rЙu<�O���ɘ}	a}E�]�B�׼���pS.�_����
 RVΆ�u�?�oڿ`J`P��e&��6��W'�՞��4��
+���z/�!ꎵ{I���̚��s�M��m��pϹG>�u���P��>d!��-I���$#& 례�_K�fm!8a��U��_�����Ǩ��L���&���>�
s�������6°t)��r��m��4�I�#�;:�c:t={�P^��7`����C���=��a6^���x��(@Ei��#�=�b�Ee@)Ax�樬E-�� �8���t��!�+ޕ�޾Q�vAF��;2��d�Mq������9�68
�^��H|��x�4�ps���3Y%:��X��52�?� ^+r�����i�;�v��/iA�]�3�ˌ�8 �"�11Kp����c������n���U�"*�<�k /;w�z���x�z������7��X� �y���%��괹ޔ��4�/#�	��
�����^ �"<:���Zu!^Ѹ'y�c�P�Ү�j���es��ţ5�����^��`���eQ�5B=�7��Lhx�T��ﮗ�~O�  ��f�<����5�+�� ��o..�du��">X/����x�A�r`�9������]m��F�?S��1��l�L�UYo����^�u{4�+Ȭ�U?T!B�+L����� ������s5,]�Ԝ�^J�08�m!��*쁸CEۜ��+*ƪ�M��(��b�X�b���u�)�͵^-�x8�9�x�����������d9�}(Y"���E&�ʐ�p� Y��s�G�oQ��*M×af
�"�zPt:�J��n�����ymYc;�|������x�1�"ۅN{T[w$����_�9�;�1��:Aи��;�S?����t�kO(p:@�����U<Hi[�g���"1G짘�)U�
*�]*�/;�ڢ��3�2����rR|:T��k��|���s,^�R�䣰y�g^k�BAj֯l�)�5��~����͖6<<I\���in�/���\��sG�*��C�׎Ӫ�&2n9ɮ��J����޺dv��x�h��{�@��GB��{>�k��Y3���x�p]
W��+�7�~H�a<S�s�+��>��K���	,k%V$��l"{��+@-|�q.V"1Rv��E��h|��y;�7{*��ؔ<�Txp���wL���A����Dx��l���=�@�)��HI,�.��Ъ�� D��p!�(C���s�f2'��̂4��!�� eF��ؙ�7Xb�W�SW��ڎ8c�B�� ,�����7�S����;�T��+rNsȟ<�[�#��Gю�<v��S:i�11.����7@�Q���n�&-z�S��r+�B=����]�3.�q�F[�h�-�L�̎�U����u��Rڄ�ޔ���t���ɄʵK��4n��/�����.n�8�ݝc�E�-"�_x�)�f�GԒ�
�xZ5�eB/����I�*or��t����ZԠ$~ �(r=̂H%��x�Ppz˱y���`����7�œ����n�5��� W�`���k�'��u���:�KB+U+��o�ydÀ-51�.�{k��{��q#��
��R�����G�Y]�X(y�.ֱ�>2��?��l���������ך/��,�iZ��OU)���RF��V(��C�A�n���b���&w��)�
!���B��*4u�Jjg�� ���L������v�#�b���_1��0�2�!�9.1lX����5bҦx@�%n�#���볣Ԅ}��=ϰ7��# �Q�	13��^�Dy���[�湠�o�7�`o�C�c���Đ�1��Z�g
��<�U��%��
�8oC��P$C ̎�A����V}�;��3�ؔg��B<��8d��ih����74���!���LX ���b�r�-���� �D��P�3Z��hT7�
�x�<��w�7JiV0��k��	�w�4����+�T��b^�zBy���$�	�z�xdPʸ:J�y����-�<n�,�֊mq���N� X�R������u��x{O��ӎ>x����$����m}��2C�^K�����]0��a��H�2]h鏈t�jm�O%����U^7teG�y/s�F��o�5�n�ӒŲ�9���J��w����g ��f��+��Qp�zwbb��3|�C�p{���w�-�V���$Ƀ����·d���5�ngN��Qvf�%1p�8a�Gk�b������{��o~R-�h�8Q���]7��=�ܓ�o�芚7�t��A�����/�?Ñ%[ڄH�������1M��ٟ�k�+���o8����Yrs5�d%�D4m�(�K����?S�
�("Ő�Na<w��|���QUoX~wS���p^Jo�ϫ�K����R0���9T���N���82�e$g��򠙻X��xЩ$���"��B}c���������T)׀2 �X"ȥ��ݡ���=q����ݔ`�����ONC����y������j�{���Iu����ɷ2�ڹ�&��ƴ��`9N�Q�,\���nةA*���N���	����0dۜJ�-&c�~YFL��C&i7��}�/\6s>[�ACKWy�ɷ�dy�qT���n�K���/����4��M��6BH���'>�h��6x�-��p�۲ɮ0Kuf�2:��s��B��b��>�u~0�,��U�t�_!r���I�������IƦ�O�-_A"�|�TD7���c�]P�<�A4���@�k����	'��>�Q�>�~��m��[F��7�]�ŗ����ŢBs�}��,�ӻ�	��l��"c3;t%��CRl�=�P>�pd��ZpMl�y^��Z$��>hcR2�@E�8�	��1E�%*�� szט������dr/�+ף��1��Ǘ���_������A+��Qb����-���H���TB<���ھ�
w��cv(/�Vյ@jva��_��n��ĩ�0J��w[i y9��P���ܘ�Ÿũt&�$Y��cSE[B'*;6Ƅ��'ֿ�޵���;uu�D�v0�}k�f�f.�jpP�V�,7M�n?�4�$����'N�#�5����DF��� ��kK:5́v2豯`9��l1gux� �X�������U@װ�+9����3|�;�q����7���Z0��0�|�8�(��&��=W΀�R��=�S��BG��2�� 7$�e��H�?;�(7�Ӧ�e��a,�ޛ��}~ۆaOY��*#��&'��=�D;�C��9):ǬZ\�n����E�k��6�f�.\��.7�ͳ2���Zn�`M$j3���S֮��lx�|	C�9
V2�W�`�K]�:9>z����H��m8-R��;!C��B2 ݚr3n��wd�A?_�0$�����TPg�Ď�n}ߩ}n	 �z�k������q��5:�O���Qc@MfҢ��J|*`n��*,s�5f��q^���@�������ͣ=Y��roi���!]��܂7G��!�y/d��(���SD)E��F+�'v��-�e� &Hx�Q�v.���;;VJ��Xm�:[|O/�.(�����!�xC�\/���3W�<���I*�䥆�h�fk���������/l�Y/��W���G87K&,��򫅺����n|�υ��]������L��u�R��U��rf�o�l��%�7��˷~o�?�c�����Xh�"�F�M�]�^��7�J��E��"�"rc�����)��D+WB���IlP� @d7��(=��ID�����ś��9 ��iEǂ(VI@��z�}��J}Ҙ*���b�n)�tn�Z�2GY���Sf��9�D�E@#4O��� 	��Q���V|�@�ҙY����<��^����zn�x<^��w�ұi2mK��e�(���j��~�������ŴÆZ������K6���X7j%�y/���S+#��sxe�!뚝�l!2�)<�-�~����� ��-����fߋ@D�Dأ_��i�[v:6E�(�;�%��[]ʗ?졧	���%L[hM1j�!�i:���㼊�	q�O���O��bL�LD�e��R
�mG-&���꧜i������r(�'p����<7E^>I�wЇlLɐ��Z�z���D����=6��`
M��^z�C3~�[߾�W!�f 
S�I��{~�s׼ �2������[fT%���ܓ�myQYA<�ѕ^.���xQR��s%���`ъ_s(=��B����&~�a'�"Q�{x����TkYw���Ce�&;>����!f�˥
[�`������SI%�r[�*vc}��jG8b-��[�.j�p�9�.w���M(�c�W�֞J��~�h��r�|$���7a�	��&e��|�[�W�٥������D�~���p*���`�KQ���:�l���y���hИNhw5K��:Y��Ɗ��L�*N����g�����C��U	MGc�+Y>�ej�)h��!��(b���9���j�l~ʡ]���T��1r���q��v6�E#�o�i�< 堣0��H�������d�q~5&h��A-`��^T|_��/�U%�L�7B��c�&�Ro0ₙP���V��=EY4�vH��������Y�t�3)�[��wER{�	��;t��%����HLk�m ��]o��Ýꘜ ��nL�R�A&90 �����1��V�T'N11@;3W,�lNլC�R����s��8d�#9G��t����@�j�� ⭖P�?/�V����n�R�����b�H�-'u��.�IB�b�n"]Y<�j_oh�����' g����)�� v�iKR£:~�I�)GU�;+�B�Ҡ��Ccc������WoB��.A�P�tx�� pV<yb���ԝ!��cygܥ��-��?�Q�p���Į��%8z*�U���c7��$ŏ�Z�0��/�B��4!; �"w�΁�|���2���{h� �kf�K� ��W<̾�i?��QlG"~Tc��uX�$O�f���#bm";>��lX��Ud�OY�,-�/k���*�2	9����!���[	�WT.i��F��c�
��K�c�d^�-~���y������uP��\��P�\|�bu��yәϲ�����I6��B��P:�~ Ǒ�h|g���%i�S���iL̗�+��_�ڦ���b��"w��n$�R뼕O;��zۣ��SD��S�I�<2t�} mRe��]�|?�nJ�ᗈ��"5��~LD���	C|aO�7�>q6G<��	��a�2M��
ح%��Pi� k�*"��3���q�=���WҤ�:��G䔅�y�H)�z�f�gPII��v�`�k�Prr�T��2��������>$�s�Cf&�2�g�ۛ�d�TN��1���hr1PR5k��y�kkm3����y�.�=�Bj���jI[��H�Z�O^
��0�
�j��G��c~ܘH�	��>,|� �n��.�����DW�S��2�0F��&���<.
���ϼ�2���/۵��i!���#������aZy@��ķ����ғcTC�o�s4�ʙhN����X�O�b9�z��m�����5���k5}Tn3Vamh��N78�9��͂uW�p8�����K�=���\���YM~ݬ�,m��_�0�aĞ��b"��$��fYH�>nM��6��x���h��( ��s��ޑ��ݩ*XKmY��A��j'(L+*QU��h������(U��`B��N	��n�%p��V�K��G�����bY�`�t Lhp�D��le��X§Մ��+���OJ�I�Z8�[��W�
dL�Lu�ƖH�k_C��r�#�$f�&������2�H:攻��Z������>'�Zꩊ��^�obb�T��	��m篊qw2�C '~:� �ŵ���w���ٌy a�^��0�>.<�y=b��<r�hR~3�a��e�
��� �9f���ؘA��l�#���L�t�2���_6��L�nRF~�I��T�7��l�<m�)�<�е�t[�:�ПoZ�7?�DVXBMF�$g? h��O*��Vd+��*>�q($�;2���+�Q/G���8>�S0���.����^�V�!���Xc�x )��p@�HA�A�feH���� ����﹡�D|��k�Uk�A��5~?�OF����B��%�tZ�%�/SD�����D��|�o�>۩�O�ܱ�x�k�%�33��^I��뙺6��x�f�ΩGBFe�e���t�i \IQ�����x� ����iӋE����ӊj����u2��3���Yi�����qa;"��lh��0�M-�@xi���쥭�&ѫ��=�U��.h��3jY�� ���ؖ��ȟ>�·��I[�6�n��F)�>��2s�~��1�Jav~��S�E��C�7\�Ϙ&��t�a��?n�ޥ�]���57AVI����}�&�Ķ�C#d���e����|�p��H���Z�ֵdI��!b�`�����_$#M� �U�GG��Z��#����]�H�M�NIb�Y
}%e�U�D�h}%.��4E=�5�!��JNi��B�>�#\9�G������>�J��5�/3�U�ǒ@��#�U����/'�N9�.C�Gj.�6��|R��Sa�
$Iޔ
ݏ�"&m	[)���
�x�
�VH$�t��O���D�ٞ�T�Y^g`CI�0u:�UE`�`��	�=}�
M������R�t�-��v��@�;Ne`x#dͲ�,"��܀څ����?�:'�����)�zo{��3C���G�8G>�H?��(�/�,��P	�^N�nA?޻�H2qw������ܴ�޺=�!��E#R��G�Z����\߲u���~��~"�ʺ&(s��h����N��$���d�2��DR�4&ٲVc���0\m��x7��'��7��J�
��v�(^)�^��q!�6�ݩ�/���Q@>4ZF�� M��@S �q1�K�����A^�k+����Ej�m�5����0f?��5tJ�X(�<͜1��(]�<�y#9~騤���������8�:P����_#�ϭ���b��[�"�{�W�p<�]'X-e��;��B�����#��4%�v��Y��dވ}/0KE��]��x� ��n�2���0���o��2�z���a��G�:��>�X,��u+�l�R�2�����r�.�F��qv���4��Vݢ���Q�|{��p��Z�h�P���Lq��@T�?���o���V[��H����%��Y��������F7k��2�5m8��\�z�ɂCWI�a�D��y�(��c����K����d�i�M�D�g**����W\��.�}^׼��D�U,�1tԼ٢z���O����lk���T3����N!q�1�����6�-��`�2�j-��u�g4q���	.!I5I����LF��/�$a�\�W�Mn���~�:(��3���Da��]���X��������X2T��#D��sTB��]f
\c��_�~뮚Bn�ݾ��Q��#��Q�7F��X���B���N�C|[!kR�����J���[W^e��*2L���N��M��?���R�̨psv�-j���E����ﶁ��X��P��[H|��Y-�1�i��B>9'���Ƌ���Z��{�~�SՊt����,�O��Ճ� ���P� vJb��l��Hr H�a�Ӥ%C8�G��&����Or!(u����tN ���)��H�{�^4������*�U !S�-y� 6�=3|K�T���AQ8J^Xh�6����F2�S�m��>G�Ƈ�9��ܽ�C�j��k8�Q�U��Q� ��)�O�ˈA��d�I���S"Mm�2ׄ�;A:c�[(\'Z��j�+z �v�_��GϹW/�� ���_�\�R�$��$=�r�����Ed���pP�{�A����	�'z������+�Js��a��3��MBw��i)��n[����C�A�z�D,�Q�0"n�y�S�e_=�}Lt�'A-�m뺶$f5/0W,1A�~����^�;Дշl�&������ܩ7R:;�t�C&6��Oe�c�����߀Q��6Oʶ�L�kI���$��Y�:�F�նl��������$�1�Y'�`�覺�m��.��f�"p��hc̠��ꎧ`Ц�J�c��&XJl̺��J���f�����0ƿ���NN}�rì��ݱ2�?�u6��
�P��b����/P)e��?�NZ��y�b� ���qq�%�rR=�����Y`�Y��p�&��7Зt�_Rh|���mPC�j��*��	��&���|��|O�1R������/�a��������ƹc��Dx1������>����y��X�<�9%��}�ۉ/om5d?*j�y/D(T�_���ULx����my�[�\��)x'a���A�1���x�>�wXC�j�y0P����T�MѵJ���D�Y��=�׷�F�֣Ԍh�^�1g^(��'�6��XˀC�_Z]�'1?;��`f�����
,�x��S0y��l���h��Z���O�Bf�ߕ��]9��%VA�L�cQQ��@��}��犠q},���ڕ y���cv"�g�e9L̸k���٠ź3�YE�dե����=mم�}����;���ل��:Ȩf���XZS�*ā�����Z��<k���w��t�0�!�� ���j�^�>〨����GA%�{��x��+��+����R4��J���[����xo���3� ���VN�"�c�f�b���������ˈȼȽ�So9 ���M�Ө���Qy�IJ���7���q�Oe[أ|�BQ����y���)ktq��t.��w ʫ������	֞�9n��.��~�)Q_b�LZ�AS<I�37�o�A���۠�]��J�9��;>ʙ�V%C���V�m ��/�"�"׿'!���������1�@b7?�������4��
�_���J$�i0S�gI��J�t�xf�i8Aμ�!!�_�%l�F�lΝ¥��/�*�sw�	[��=�����"�@�ZX�	���ޟ*2�ZU��=|Y����m���.�9^�����L��Hx��bG��ߧ��хn�<Lfg��Qv���	L
 Ʈ�u���[����H�1�Ӏ��zΜ��1
�:a��/l�<�D����������u��yU���K�ڍ+&q��?�ՑP�G�̹�(o~�u���%`��=��Ub�fm�|�X$W�x�^L�%�U��En?Mo���38��=�Y�K��}{%����C�dP��;UdKEҜ�	��UȺ%j�_���sXs���y�~�;��P��SsnJ{eX,��G֋\b �������ǭ-���i�+��~��0GL_��WSlZ�4�/͸yw�.�vº��.�ߢ��K�`'R�mb�� �8���I�����8�P��< �����՘v��u�\�JPB���1���rP�۳�Ι��728��>�Pu����	��=����V����H�A{>cQ;@#La8I1�T�����I�P
��_e�r'�{n�"��{	��~��}:��מ&m������m7���եc�k�����5��媘� �%������u�c���	�APý٧� k֧�҇�%_O3K��ˡE�@@�*��|��a�g�n�Q��q��%U��JӴ]���xi�l��E"A��_��s\[���q���a1�F�X�!���t�Ny��ʥ>mFj�6:�U����b�KF�x�(�_qz�����rS�!Mp�5�U�R�S��Ļ�����ft&?f7af�	Ѯo.6��3jٱ��w����Q�_�;�=,��	�Uׅ�,a�Dt���z��۵-�ƓPh"k��:4����u|�1�X�!��&s�K:����mQ�>����r������#�fل~��C����C_�y�$G+�I�0��H~�CQ�g.��D!���	��,g�44*��0w��Y)M�m��ZOb�yt�fz�o[6R�(��=����y��S0)�c��`F֗3�V6]�!1<�C˨��9���4�W|�q���̅�ޏҝn����#�t���[d�'"����U	 ��PZ_a�1�,�DULA�ި���6�)t�B$܏��	�~��(��%�alo����a��1(b3�>1>�[_{���7�a��(������ح]�����~��4�!���je��@.D��nWVW����p�4 ����+aV����s��׳PE8�ز>��wD���A5����g~o�3���)���p:!^���y������!X:P�E���]�c6?Q��z�Jx̆�Z3[�Q�pA��.��g��� VYq�Dd�\ ���:/�=���1SkZ
��N'"ݶ���$c�b�%�"��#X���f��r�LF����M��i�m��v�!�O�^國|;�+�ʤA�S;,�Ќ+|��G�7�74��/��ԕ��\]8�l��=�p	��;A��_���pǞ��T�� EO���
�(bMN ��В���9�4<�������=��Vj���s�ɵ�x���a������Qo"��!�_~V���̥a!�ne}��z����E�8�<��^����w]J[!��v%��|W�z�%���)7�;!��Ԑ��X���=��EQ��a�(ƾ�������m���`X���nf U�;��Y�ү(�f�:#��w(%�${oFj�~�9"���D\K�n�a�j 	~�a��߽yi{��]�\��]��0�h��^��6pB54�۵�BZ�A�)V�&6�U5��I��5��Iݻ����0'n��wk�����,$�
ҏ60����
�@|�x�$+ ߐB��1崊�,�*9����yj^d���;�N�g��K���g���_}Yc��2k_ˬw�́���d =����l�z�f�r�<�q�7���9w��$y2��<T�䶛��H=A�c �K�J&���`u1�{r�����Fl��(�H��h/W�����v�n�%�
��"�x���͢�����`�Bt?-��1"����^�����K�ϛ�$��^h�:@w��6��89
�ꉠ��֞���dz@�ɰD4�7G����x!V����������%��m��!X�x�5��I��w��֏,m�L��X�����ϛ�+ ���Ѵ�8;{�5�'?�>r$w���c�o3�^[58q�I4e{�@��vqe�6�) �-I��/l���Li܃�S��ᖀ���"F�gΜ}�q�X ��(I��]e'\�nI �Q��.����NH+�H���FEK�S�q�� ��vW�K�gAԀ���C0�EQ�*2i�ԷS�W���ޣ����9X����f�s�]πu�^��BR$S��T�=ҫ
/�drs���lt2����&��s��`��5�ԇI�����%c����w�W�l$�I�a�����Y�LU��k3 m<mn�Mt���kY�5o9<a�.��a"���B�f�T����л��xP�NQ���g��HD[y@��At�AYz���&2�w����ᣏ��[����'��R�9u��5��dX���Չ�1���F���U�{��瘁6�K6M.e�3���t��\ "��|c�@�؀�z&��0p)�j:�~Z�y4�c�ݺ��Z�)�ۯȾ�+��%�x�֯��@ 5�j@�c�&F�]������S4��x�y�U�_�fY�^zjҘ:�Ȟ8�M�����I�q= �$ק��TJ��^���*�	���O~��O qTꖃ�ŷ���r��{,�#�	+Υ�ѸI������Zu����M�N@�����x �kjus��򾑵��yD^���d����GͿ�qw\Jւ.P�wc��� ����-"�,-u2�v��X���)�ќ�49\~�N�u�=��]Z&lOu)�����V����Ȃ�31�����Οik�,��/��__���a����7}�`�>6n�����'��w�W�u�,���s����	�=���!iOn;� X���I�K�I��;\G�f�+gK�"p���"%zy����XټzY
��l�)l�y���Fȳ�����
�6��تE��L���m�~�#q@���>}�����ƠlJ@<0uH�:��ׯ���M���
g솒�a�d*Bܔ��Y��lY����Rk�k�W����r���jG� '�5�0;$˓��=]�Τ¼O�kK��Q�� ��b�p�3�3Ⱦ׮~2���D�%�ώ�G�j8V� #es�Ϲe�O|\�4�x�͵�IP����"���U"sټ��G�PenJ�Q�|��n�.N��?�jO{@�x���&��O���Q����cd��;0�#G��8��<��p�b:��}L���%D�G-p?ّJ�n=?�U�}�r����ڬl}?C*�3 "���E6��!�C">F�@W8���Jŕ8`y��c���*Chk����.^(_�3M�Ž��ɰ���I~g,�A
�a�.48f�;\�94�׸���#����T����/RB���v�]���ϫ:�ϫ�Z�:�Z`��K���2���v���pi���j�"�O�c�Gk��h(ό	>S}
uCYk�H�^������=�����s���'�B<T5��ګ�s�Xr3e0���;������|��N_���xW�Ϙ}��!:,N6].��ꖸ#5�rS��haY�X��E7���s���A��ZL�lr7;q������HBg;�B���y�%{�Q���:o/�qTO�!���ƫ�K�b�z�U**@�B�[�~}�����.3�b�QN���/�����P�<���۸�)k?�V[B&��#�<��	�VT���R����̹�A �Q�J4����{��g���;�R��tKV������ku�"�tӓ��h4=$�j+��xDװ�q�@�;]� ��M����ϒ�5�9�0q�.���΄�H4�#*��֞� ��_�^/�Q�,����D7��K����������8!�Ο�r}� ^��9��.���q�X3**��v����l�Fw]���v]���c��-
�nT�i��`�\��>(��Eɱ~m� :����1[��&�e�HF:�#d��}�]�_����gTסL�O'm^��xK��U�y�f̈�[� 6�{��󫶷�U���3�a�|�E�
��L�¡�7o'��>���OU"i*��K@o�4�����o?���4����3ϐ�Td���g�ߐ�w�ۉ������U�A,�D}�R+ K����'�gF��V���
�(S�9�t������>tR�j�+����O������S�	a�*&ض2Y�틟�T6!�`S�H�W]pn�k�N[X\�k�Z�������x�nydQ�xȑ/1�9W�tD��7��Ϟ?<�/�N�"�KYk��S����W�C6-zl�r�q�gIs����+k�[؛O�5`5B�qk�u �կ�&�D��(0o�X�����`ja�Q-]���`�&/�~ƎBNb���sB�Hl���pI؅��2����)����D��XK��n��ݦMʣ4ų�)�@��4$uV���4�1�;xo1���ln�.̾��>S��-.��t��&$�5��,�������$I�ƣ��}�vz��nь4���Q����t��B��L6F��]��m���k�#�Sl��jCUe�u����$̬vJd�-���@3��*��;�B��g����~���:J��-t�#ε��C`��AL}�:�ڝ�¿R麇�:,�⌃�ۖla�������#�ev-
n`N��� 4���3�_A�n���7��?��pF[�ģ��R�j���D�.���Y/�n���e���`ZZ���Fi�=p�?����j�����1D����;�V�$Dά �w�d�H�BJ$T�"�G���g���|��?�S|a$�G�j1^��s�	�O�	�$�&R��1ؔ:=��6�9 Y�UoUC䤮�[���<��QQ��
�~��|���_W��k%:�o&�^�W޸�p(�`K���o�����E��lR�{�]%�xR2�r5�_��>	��Š��:����:�D0��1�&h
|R8�J��ӯ'��zqp{����!;��u���#��HS��Q+y�D�ո���\J�х�%��h����w���<S�40�腎ӹ�Э�<k#
'dJ�O��(#̚��q��5I���gӂa�YQ�=I����
{_%�*����;r�
*��C��;�pNc6�n��0`6u�.8"���:���#�&�Yj`�U#f7����T,�p�����7$�i���Tuyk�,҃[_q�۳ǣ�����Q�gv0�����M�`�[���Ys8��0����eD�m!��;��5�3���`&ˉ�k�4����)h��qjx���ާm s2:^q��v���q@
�3����H�Su�?�����_�{	���)BW	�(bQٌ�С�����oB�
��e�kϴ2|-��[�}��`��C��%���[#	�K������0�+���0	��\U���>%�ZBc��G	7Jq$�;Z�o,r�BC�� ���w��PA�Vuok+o�&��Ł�v I^B�yG���r7W%1���53����#���b�W���ǋ��n�ި���ꎜ���V���'F��tX�����	�Z��°+��ň��2���l;��OX��f.�;�_#�]
���)��rɞqf^��@�q��7P�0��Em�����#��˓4��L�ZP�����-��x��6����*�'���j:a�/Y0�Br���C�2�~���Zm�� ��?�ץ7
⸂�r���6��0�~��C.e�Ee���I ��0��	��_�̦B���nO/v)�6n�B��Vp�:�+���x�_6-����i��"k g��̎]�«3f�c~:8���~� ���@�o$�劌
r 3�`xh�b����*w��B�`�M������~9׀�I
�#k�!k�ܸ���?L�xx{N;e�юѳ����v%8��D�;�-� g����X^9~q���S6�u����S(�ү�����|)��	�\���
����m��kl�p?<���q���.ƚj,�p�[Jx5�ԥ"��$�-,����E����'��KG�[a��涭<3���k8���ۂ�c��*K(��+�������w��q��v�
��:�Q�Ua吩E1/6�W��Ƒ�%������g���V����ӳ��5��X?1Q$#6���:�[���@��Q|�s���ʁ�-G ���?��[��x��R�ٳ���6ԓ/`6T����Pw�"M�~���XE��פ�/�#tF��Kף�D�Xo׍�!x���q!nT���`&[?)k�k%���o9j�G~��Q�C.����"�Tq��C�T2��ՇB���U�7�)����@�ݸL����m2�t@�d-="�,K��A�¼�Y���ߑAml���X�a�7Ou>��V���89r*�B�C��#�KU.N�4D"���I�X�G�l-&K!���'VX����R�fU��10�W�b�9�m̊��3�뤓瞦 �)n"I�����]��:k���GPDoӳ��F�@�d4�����:�؅m�ԭ�k�����iD�x��WY�tK���x5[LVrBŎxY��{d�bf�������^�J
xVu�!���k;�Ȧ)EoG�+iR�&�p)X�vzϑ����J���M�69	�w�^!6��R˫n�:uz�]Zb���I��m������6l(�nr#�����e�R N �K��K¸��)���ՋT���̟������s��9�����dc�����?��1��b����̭���W��ܫ�`�n��X�%���O�._.���ӟ`�@���ip�UL�[ϫ.<��"q�HJ�g�1���W(���{'D�ו�ŧ��K�IY�!.{�@����p�R)Tc�J$���f1��s�����q�=g��4A�Y��!l��o�)�m�ks���]l��;]���'�e^�B�G#�W��C��.v�Q��Z�I������D�\�X!ҷ=�{���E�T6��\8�Z\�5$gY[�匄�`�<��EK��w�OE{����\��8ó`z�����@U�SZ�E� ���y5-NV�u}_���`��u�UMA��
i�\��K��2/��1���a|�OZ�Y0��]�Z�Y"����G�W3��vo�|Qwg� �BB���*X��~��ME���c��f�g�4����3��t)MK�������p�P�4d�}�1X�i�:U��E�+��I��Q~	.����;���V�~���.��%�G��>v��@JAĐ�E	@��:K��"o�`(Jh��t����e:n��ua�S��B���C��܈�@�c���{�g�0WP��PaS��5 5�XX��/m \���""(�m<iy���G�'C=jz#�n��f���M���1�z�-e��~�=�Y-|�re�G?
�9�%|S�O�M����3j���2_i����Cň����5���H�5�`6�V>��@�ELǤ=��O�Ev��4=��bI�UP��K[�����EK3���8�J���Ւu��/Ғq��c�ۋ�*N�p��V��;@E�s�{X�y��y���^h�C�u�(���J�T�$�n���N�y|A�!��+�-�˾_��ͭ�ݧ���0��[������7Pp"���y�`r��]�u�mſ��/5�,5>��X ~��:�N̳�#S�:w6�B�L�M�@�3�]i��-�h)`�Yߊ��"�g� \�z�S�<I�����4�[��⍚r���_�K�
�ڍ >Ɋ��D5����|&�|�B����i^h�m���s�jF��bEܯ������!o�m��Cm�@�s���'����ԛf5W@�����@I���:q<�j�)1�l��M���}V�ӏ�����
�,�$�:��5�����7"�H��@��ua��:��k�s��E��:�[�s,��Y�92����/J��̵8��"cG;Bf��2(�>��)�g�D?)�>U��i7!%����g�w����X�qr�#�	1��au��86�ٔ���1��mcg�׆�i�+���^BJ�v�71����^�{dՂ�[�h�]@����} �t�di̦��9�g>�z�F��SL���
��ҭkSϱC*MNG_w����D=���֦�w�5d�ҷa&^5��H۔0��b,�k�g�#gҶ#�`��Ǚ��K/팒]��0�	�����R����\gP����0�C�=�IF����i�u-5t�՗ZeHɖMе��2���OӇI0_��-�Ү��Ŷ�;���ڞ|1,�9������-�g�
]�c��]�%��K-��#�1j��]8�D�8˭
�mKC���޴�������FTȡx�>��9I	r/��d
��i�W��Nl䈆��X�xH㎿������� �7��Q�m�T.P���
k�,�rޯ���,��́��l��[��M��&��b��=��~�J��X-�K	�A��^� ~KHT��5|��XE�W:�[#�E�ٹ��`ph�N7�"�7t�I�v Nj��Smb{Nk#b_�S�5S>k�����s;�$Z�f�`����	�埯��S� ��Clzƒ߻[һ\������A7.E�%�m`ߋs�:\�8������ҩ��5=��/!]��y"դmස��o�nö4/ �᪞_����c�[��o  ���jcv�79��c&��KP����_�F��D�(��F�Z;Z~à}��*:��=�-�|��4�p�At���zu�B�_���Ǔyo� ?�ȷ�,QE�I_?����[+��Ra���(�#߳T=�g�2�#��tE�/�$25v��,ۈ{�ִ�Y/dS��۾6��� N�����L)�$I��,XB��$V��[�� �L�0i/�v��Z��D�t��6Vې�%��(�@�T�g�ы��
����c�N� D��>$}�+��e�Kz�9W]�Dtգ���|sm]��u�,�Y��o�vc�ؤM�L�9Д2��!?��6��ΩF��6v��}�T�m����lC
V/d����w6�t\cf]���R'��1�3|��Qc�'T���2V����`v�xD.-��Pk�P����Kw7;� 3�J_��+��b23a��Q�5Ƞ���Ҽ�I���`����#
�(��D~��o~�w� ���/���P�{",��ق�wdv�[<(|���pUݚ�XQ��Y<{��3LSlt����|m��]{�Ү4Ѓ��}MAz��y����bHt-b��f����_�r��I{r�� ����R����ʻ���]Irb�m�w	F#)p�>B�'��0{d�f*��u��}ZM�	r����!���`ݸ_�2��^���qxLrN��,��\u��2���R��#���?
�d������ʘ;���x'nP��s��n<ד������	J�ε.���(���h���V��9<��m�K�cVC��%�
�0�j~��`�l�xQ�b�s���v,���XA����r�g@��h�:4��x"lG�X� ���դe\�߂�?����>��F�=�)ԩQ�ڝ?�O�S�#�Y֥�1�^��O*��1.Ⱥ���̀�?��E����^��`�io�q�����G�_ Or�VHm����
�@/�?�<��-���2�O�=±��Kp�gP�X4���P1=
s�IIؼ,,3j��`z7�.*��Ξ^��L��>4���9��y&�f���$���p�x����ͼUx��9�䌬��q�[��-�Ýے�K������`/%� �-�s䃃�<C�cr¯ƽ]&�V���)�M�+d�(�sG��*�����Yi��"+�|g�;ۅ	c�pU
�ʖ:��_�|'a�����?�_�Z �X������+�2��W��]�)�2{@Re�&*��?1�XN���5wu����XLɘ�ifx�%��7U��}B�&���bn��Mؠ��PY9��@��T��9�JO�_��r�jl>r��A��v(k�m��V��Է�ʝi�@�Z*�NDW]ԭ=]��hl�ھL�USO�T�b�L�6���ؙ�!SD��?s������|Lv��7�/UЦy5���V)�8�8��生��\&-�d�)�r;�V�qޗ�i@�AfZôsӅ�T�(��u��c������z*f {Ʈ(�GA���&�[�=�`�J�R/0�T��@�����8�|��w��L3��L����b�} ���=���J�f���Vǋ~�X���7�ź*̈�n�"Wv�ok�<�E�p���6��x!�Aɣ����ߙ���	F/a#4�ObV�,��ۑ��W�T�+�0U��1������N���q�1�[�ȇ�>�^��!b�6�o�0 {��,=�N�r�מT)x�;W�dĆ �i����u����}��}c�A�%���˟��ح�L��L�`=�/��|}�'�g�W�m���'@��-��xHѪM��6�u��cbؓ溪�)�	�8i�o�/�]~@��W��5�"�%�RՒ���ѦE(++H�WCE*��R~&��~5�h�S+�z�ԍ�Ce�*��
T1�E1�t��>��,4[�az$>�7�/c�d�����M\�OvRvA��ce�y�U��{%�ڋ�A�\-q�ZR��8�z(�4 �L+�Hn�Lv�R����!��N�MH��b3�)T������q�q�%z�sװ�Yy6���v��W���Z{i�G!�<?�a$B�"�fM�N�!%!���X�ʎ��^�E�|
���6ÙJe���25�Ph�俲�����<���	d���7<vo:��9ܷ�@���ށږ ����Ewr#�V��~�^����_7f�M{52L�bvE�����`y��������얔һ#Ж�ӯ+����I�}�[��V�J�H�P*�)�_MCG��lp!���[ДL��x�$����nr���B`�^��u��ͷ�c�'Q��9��[�lqW��+5~tY�00�u��*�pD�Q�Ly�h�T^��8:�b�ZK5�U��潠�e�`Q��."�|K���,t!�:�nh�v�`�A�F�!-�>����;56Q�֕�0���U�^����4�_Zb�A3��]�6m�\�䯣DD[�2,
��Ō9���$V(Cv^�0�|��7����L�ъ�%��9��I�����k����9Q��~Z��|��G����|�lD$
Y�d(k-9�ɘz�幧�U�_{U3��\=�]�u/�|�ǎ&�❡3I�=B1 �Z�229fA����#���%/����{��C�X5)©4=iG �h�3�OX$)7pqQ�;���`]{�J=���Y6�e��Q-n�K�5o{�m��[�Z3eF�Ϧ�͇��"�l��8���1P&�G��=�o���	3L.
��F���Ɠ��_j��8NDi��U~��]%�S���*�O�Y�ޖ�T�r.���S�k���h���iB����%z0�BVMvJ�Ms>��2>
�h�8�^/�����^�K��������QJ��Z�B4�0J:2�Ua�Š������i8E�k��5�s��d�*$k�x�^��7�ȍc?��"͋R����eI�1t��	О������"�ߴWb��i:(U��~oA$�:�z	T�POJ����YjQ|7+��M���E�<��Sp%9�+cn�d��u�.\4��1N���?�^"�Eߙ��a�,�Yn�/.�$�$��#o8���
_�eU������Y��Q��Άr�C��UPc����	W[�u��<��7��ָ Id�p�"u�$�Y��zҗ[�%N	[�bɬy4�QN����~�CK1&�|j�+�Q��H2�[���m0vgE��C&�k͚JC���S��{3�Ƣ�J���U���4�i�v80�=��/��]R[���X� �nц=��g\��u�D܈��FZ͵�=�oAkK�0� �r�HĞx����)�kB��1E"]��o��D����������hix@�ӭ���W�[�{N=�&��<QgS�Ѻ�s��JcjG��M���~��,!��v)�I���-���}j�:�(��"Ia�\a5V�۰�9��ܩ��e#`�'���NpV�Pe�Wz��L.����T�B�|9��Z���"��S����c�Om&�0qvi�8������Q��m��=�>.5}�%�_�BA�%;��I���F&	���~.`]*GZ� V�xY��-���q�#/��W�:�nP����)�t�+�.tFQw��r2Z�m� �����eOH!�����/�q�<^2� ����v�"��4 ������)G��s��ǿD���!���n���u)���JS������&���6_e�G1#L��їG�}���9��ߝ"s��,����r�͎I\�ʁ*�M=1C#���jAɕdW�.�?�Y�o�f0�J��Q����O}~�V+�!��1i��jdNmG嵤�.?�Nǅ�	���,*z�E�>�֒#T�8t��T3�P&�� �9����P�� �8q��}�f8we�k������VAEP��S�W����Vb���8���8��:|m���UoqX5�����c����~��h̓�@���>���{̭�n��s	0#	s�ER�_N=��U(:#LJ\hϿ�T�,<����zb�*+�F�T���Ql�Q��S�ݳT/E-Du�MdXE��R���H�]��ي?%�q�'�f�u&�����R��bt	��Z��!S	~sI�V|���\�Y�� l������3S�4�W�Z1�b�o�*S���q摯�s} �I2۬��l���=[�F�E���ď+����Z[��<WzS�����/�#S����?Y��O�*�X�D�b���%�~�5Zu�H��U�R�(��D���N8�x��Q�AD(&5��]�����[۞?,B�/��C�~��L�M&�XK��ى�'�K�e6��3yVu��%tq��a�<��w�8լ�3�#��.��_h�mgm.���M��Y/X|EU�c�^sr���qf���K3rfG��S!`8wj�S���7p!�&�š�����	��5�P��CH���(*Q��[XoP�C�G�՞/��W����sFm=ġWIlv�"�jŉ�g�ImH��x}���\*���P��&��*#�we�����)�r������`�@�~V�q���R�R�H�=hP���~-ۏ.~�4�e�|��P���:r�����v��CQ�J��L��=�'"����y8�p�Pt���ݘ�?��~�iKq��qd
�bʅ��SC����a�	���Q��l��Ƥnܥ��e�����= �p/�	yHl��j�06E�dW/+��l�����*�T?���4+��g����#j̬�tg�Ԁ�)}IY��B/��yb溎F�K��[� 2(�5Szİ�����0c���s�o���
��H�*��۹�2��	��c�g�JL���&�5V6�^�}˽�~(�(e��"�o�����YGa��C�tܿb���,�,���$�����;�+��>oՀ�3�"�e'��Ʀ��)@=�YJ�%@�PJ��G�X�C8L�?����to�N���P���������؆nL�� �845�mk}�O�����[l����IHLIuG$�c��d���U�&u
�Z0��1Ē��qB��sR/0��q��W�����o���)��A����Crv�"�#�:[d��:2������it���BR����pwm]�V��MpB� �V��*��~(���O��Bb���fŋ�"Y.���Z��^a+{]��ᑩ挸.-��%i���;O�X5��n�`��k��v����Z2fv=������.-w���l'���W���;ٴN�\�Y��K?s��>b`����E/o���`8|�sΞg�bOm��}��g��!GFZzU�֚VU�;���4�$@i��T'J�(s�2�C�p]}��~	mV�u���?_�S��=*��w��ç�,9�HB���j՜���l��򌁜cwY����޽rr��p�R�I���hN�W��al�kqA�g�1\�ХV�!_��<��-?���
�Ы0ٴz��E|4~�.��~�a�{�;�V"Y��@SI����kp'+������<�썄B㧊�%kVk ���@ ��_��E�M�t������l�d�b\g�)Z���{���q�!���n�VS���Wx�A
�D0��ܫZ�A������R�����) �l�ؘdL4�ь�����㶨\���Aq�����b�
�A�6�ҕ/�"fS�q���4t���a6}��w�OvI��Ա�A4B�̪��������&������_b�+~R�m9�zC�*��k5Ŧ&xцT6�!�;٫`��:�Ξ-2`�R���%X`6���=�Sx�pg/@��P]��˷�|�%�K�W�֕R�ve$,�������Va�;`�K���#;G���Vz�i���͂ݗ��@G�J�ERH�V��}�����\��M]�?6�@dY�W�b�ߝ=��G:��U<U|�ٻIg��k�u�A�A9���j��$�x3U�/'�-����Ih�#��s��nl'���Á��J�8#I��I��F���&#�qR��gX����
?�V0��ƛ]D�0ź[H7Y��7p*���]�j�͂�h�����2�����V�g���~gNj��7ho���+W�W6����Y'34�5�rU��&b�
\;�8`�W���u_���#.����U�?�D�2�N"a�x3P�ut3 �j`�i�e�
�sOb{N0�@�"���V[�`Q|Z!�"�����y����P�щcqM�&�JM���@��a���?���qO���@(�W�Wo��;Х0���o���TЫU6�ȵ������8(��W�Yx�X���i{�d9�.��*��}�!��O�R"�1��Y$�Mu5{�&9��H���X�@wvl�������9~��䡐L`���rڞ��9/936�fjQ?8yP9}e��9z<�/���>^�ʛc�7��qklD�9�p�aK�M��&|�1�1�֯���O4����i[�!�IIg���������ߨ�S����b,���V���>
��������1���K����|�u��fV�#��##���)c3��`�y�Rښ��o��M���e�pJh��v�� e�m�JoQj�d�P
0ZC����4����[�0&�7����^���' �\xI�x�j0xF��P��O~��2�b�F��4�B;�Y �
�<��Ʉ�t�VtF�B8�dl�l3�Igz��p���(H�*�#n@%
*�@ֿ��q����>>�� ET��Hg�g޾�*!$����T��l���iG����M�:/���t��u� d����k��o�U�(�w��|��i�K�j��J�X�fD:r��1�ڱ�ڀ
ui�r���6���R��� ��]c*g���3�K�" ���T��Ay�L���#�ـ94�X�K��`�Kldy�x�W�@wn愤�Xt'넺�!�;J�[�R��7�X+�������2=�(�J����n�܋Ï6�8�nu��t*�C?˃%D�����e�&�,~��-ra}��v��������pS�'(��()�q�_|�=���紱���OF��&�".�9�a��=��_� ҜG�Y���;W���s߄�n�s��3�gS�%/Ko���#>ؼ�I��F�\�'�iem�,;/�.��7"��m�qžv�Z.�@�`����ͣ�\1�1����/\,pNC~$���"��3�)�pӭ�4ӊ�|C
��'`fz=��_@w�N�c7[ժc�������up�<qD�_���I����q���GI��Ts�"a/�����Bp-�]#��vD��s��U�~u\�E�T8ߎ|�KW���f)��0P�ܯ!�s[FP9u����~��qد�;����UАQÚ$J�:5��+ܗ���f�r�9LǪ�tŪ��@y����@��1�
�%��;�KBD�9#�z�c�崗U�Z~C����!�[Ή��ld��1�T	,���,*7�}(�#�,�S��F�B�ȯ|�5��y� �&�tPF>~ᲈ,C^~��ܛ+S
�o� ���NȖ	�݌$u��PH����5ʬ����&IZ�_-M[+��"��h��h����p�����k�U�x��j<en�GS闠F���
��:��?Y�KJ���W��e�\[�]pN��˔C�wK5�o�2���T�'�bߘ�m��~�BW2�+)�۲];$<��-.�� = ��4'��5T�.��<�!�Ukp�;�C�|.��g$��������ɫ=E��p��6o��+{F�)]����H�N��Z�O����V%��n_���Կ�OT�KQ�MѼ�<��St���b���⦮�:n'�Y��V,��K����
�FS4`�������i�z^��!���|B+�Or�;��c&�B�[���W7f�-} ^�����F�C�%a5�G'Q�f�9�b�X�jE	���J��6Pj�m[�"P|�E�p_slEiyR���m�A�O����T�)^lo����^2R66���L���}�9o���B�N�[qF�`���XE=��zap�� �W��C�6�0��롄؝_gc��x���S��P.?L��Lu(���ײ������|�L�tm����T�v����\Ua����?���cx��+�R;v<�bP\³18�y�b|�|���1<�ƾ��Ϟ��i*w��W�U~�Ǯ�Wv�}1�y*�b&k> �-A��V84�?�(��(3��oM�0I��k�з	���1���� 
{E`�|��� <$c[t�����|�i����~��Q��p�q�B�ln�nZчP�1�9;��~&,8�(Nk�H�a�P�,}&�3��-��F�3�S�Q�~�����2�B�ذ�u��S�F�gr�h�r��8�}���,i]������	�u����-�m����5�Tz1��N��uy�o\�#c�Pt����.�w��=�1O��u5��p~�^Z�������٩G�~�׀@�
�PY'A� D���w��� ��������vPT4�ƹd�k)�k�(��:3%��@�"[�D������8�e��:�p�M�ӆ�����_�پHPʦ��v)&VK	�I ��+�C�����aԵ����G�/w�:�YKz>BՃD<,�0�/FH�o:l�s��ECsJ1�e~K�Q���ĺ�8�Dy��I�2XZ���O:�B|��il��~U4
A����=���uM۵�s0���K-F���D,�5h�ӫ�On��[q0&Ui���A�]�����I	Wb���?�s[�.��bQ ��˭b�^�萖X����F��ء�68�.�T=�$��Ǘ��N=��`E��Yo2@@��������:����}!�{$9�ovd^��U�Mĥ4�ﳌ����":ŕa�a�l�e^�ٟ����_�v~��5'�nD�:q�*dj��|�pt�^]��Wf�ҵ^�ѢǗؗ�"8���kT���04��j�j�}�rބ�T��t1�7�5�BL��]T��rn��#�zV�����6�Ӕ��$�m���}(�c�O���"�AՕ��(�H@q�F�f�1��(F&٬L�|��Ch��6�B �Hc�N n�]�v�f�0GV���g�Q-p`�_��*�S�<��(��J���x�ۖ� ]�����~�	P
�'��XL.ӌq�{���aj���B���*�R��Qc1D��3y�_�̅Q`�}��_�=BV %Y݃_5G +�WD9��@a�f� �;8D����Tn���}7��~�i������D��?��:z��a����;�T�AVMK�G��d&��f3�c�6Vz���{��8V�$�Ue�f�u���?��hV�6�Tiޥ�K�A8ᐺ(�S�#��8�P �c����9��$�k86F���X�H�/�p��@�ə��Xǥ�ٷ�#�:L?K��ߴ����@�d�'�W�p�)���>b�iJkJg�@:��[Qx�(�n�-�W$</>K�:&t�/�IM�_Uy"�:i��jm�k��"cmQ��XZGq���Z��;�w�š���T�0�Lg�����-�[�n~�_U$�Ĝ��Ŵ�g�x��67�3�GH�4�6;�=|�\�Gj�e���-��fx��FХ�0<%^�0R���5��G�K1�ة`Q4�[�G��r�P� ]�fҠ�N(]���Ѣ��86a(P�"^�cpZ��D�
@n�#�z��i��J>;�w'�L����È������^@96(93n˪١��1�U�m.��P3�r"�*��2"�����\���S�U약����t��p�3��s��TIk�*��C�_���'&}���%���h,��g*U�;ެ�ZQ���O�Rs�\�s,�9!c]hM��:u7C�D�{����_��gξ<0����ZdRX rŚ&��XJ����g0��w����W�ۗqm��.z��/�-���t�F��ڿ�5���Ja�3%�s%[Θz�z�S�>�C�O�6����c� <�����J���`�P[��u ���#�i�n'���G�6I�%��Y|����\Þ)lr�wFvNT�â�"4{��'(�'�⧇Q�m�h��e'o�-���+�:
�)0qQ}@�|�:B��ƃ�tM�褚:g��}4N�X�)@��{	��:���\�?PZ��;�G��H�b��e
{��4��3[����`�c�� �3�t���lgtgҪ��J:�L���b��⒀���9Bvꕗ;���6fJ�#/o�T<f�V$v���,&3J����&-P��|;�;W(ҳU����^F2Di�?i@�
fgX++�'$?$��]R{�*�02z�Kh�֬h�,$U���GLd�����覜��.F�/e��+8`�>���$S_6J���4"[ BDָ����3��`o6��3j��b7�V+&=Ns��H�Y�)���S����3S��lr��j*�'������y��<a2�}������H����S3m\�av�B�h�=&��<yL�.�:�{r�n��_dГQ2�[�|k��U�܎�Eady���/b�����\�X_��h�Q3Y���5��a�L�+���^��3�T\���@��ͯ��]O'�('p;�q�K;_��Hj+Q&]�y�xF=tl�µ\v�,G���(��3t���f�r���@��.[���o�W�$���.}��k�ZIw��B�rV��E�,�7�H���|�	�}��f2]��ш�7MU���<m��!����_5N� ��r��J��؎4�Y`�ôo�c���/�Z�\�p�0 T.�%*�8#�:b ���ٌ���6�0��)�k���]D� ��v�-c�p/*d�#D�D�/�)�ЎBW4;1Te#���V������̪؛���2P�\�(I*ז|��S��V� t��A�%����+<BfaO��\�2J/�7�H��İ��+�s�;�6.O)n1������I:1`���tQ���߼��C��r�2Q�v6���$�����U�GEF�2�H�����g!a��!�N��-��q�/;Êe<�=L�7�R��dcR�
@���F�����oQog��v�K�W>.�_<G��U��rg�f�N�F�=�	����S���Q��ڡ��-�����)4��y k��,6 V_��Ӷ ׻��|Ċ@N�!��$�ʙT��XU��!J��A"���?�a��!����F�n���2��ʌ��X�!��a���Ru�1������l�?A~����;W��G���n#�ø�C�0�&~��]������ؑ�t��vm ݯBfjD<�ŃiM=��I�A1���(���X	Ȁ��0�5��S���c6�S��Ҋ��v��!���<���}c��âs!�}=��)G�N��}S��U�Bt܌���VeB��}lH換I�Mj;^�h���)_�پ9_��s%0�g<u}�3�g:2u��Η_��О �W'Go�zsر���}W�K}|�imv!b�h*�;��̐+`������QC�<՘<�@���oW��Y*���c�Ff���(����!~U��q˴��U�����}s=��Z��`�J��� T��4�Ӌ�5h���`^�(����t7!�G�����m+�Y���b
��T�/�3�ͺn�����C�l<z��5
z�}��l�n�='o�CZ����5P�}��{`�0��f�\CN� 5���4R��)k����>_<���i�B�m@G;�x#P��9���M�1Ģ0�K0�i�&@���+?|H��9*;:�?K����M�H\3�����J�Wy�f��7�7���ݛ�8/��g#���؝�M�Շ��zB6I�3X�ňuB�(�_��8�oFm=��kz�����)�"��*[�h�m6��0�Ze�]��3SFrc��L�GAD�.���U�l���.Cs��]�� ��e���MQ,��4B����.��}/6A�h��f�_�B#F E�x��<�����e���˪�_yt�%s�b@�rse�mV,��Y�^���`r�����T�QB5-q-��X�D��!�r��Rg� ���䭸7��.�}�5�	��ﳢ3�Q���=���
T�!ţ�˾���Se��[P�Plx�iر|�ڥ9���s}S�8֮L<&k��W�&|B�V�ܭy>����|#:v<����i}�]h�+��[�ޱ��*�q�0��;7&i��:q���į��vN3-؋U_ϸ��8ǚ�C����wv�[�)Ö�$����I��$�a�h�Y�2d��D�Ҽ�]Jp�I��71��;(������bm1��ZT��_��wݒ~;[E��;��sݘ�?�!B�l1�̛fTXӯY�t�a+�9��ՠ���w���Q�m��緄��N��P��X��*� �GN/JB#}���dR�]�v@P��%rC�K��e�t�{*տ[�I�@|���*��c�G�pL;���U�-��n�D���	��N��j�y�E���?�t���=��b���8JR�%�z'*�3	*MA�)c9��%L�kh�#QV����Ppp�C^\��a��I��gC��cE���]��͕�)�Xi�e�eC��a�Su�*Q_��r�`9Ǻ�֑��I����.
_���cJ1�,}e��{�T�r��;��9k���i���i1�)=�G�| ���a���Dy�՝;�r�G~�;�Tn�ɀuY�>�N�~���\�#�Ƣ��D-�ʱ婞��}�!���=��h�>l�Ӱ�SP�G�!%�(������ن��~��C�{M�F��Ü,u���B\����s���LM�+1��p���H�46��$�����֕�_��{OZ�i6o�nv,"(��Y���/�7g���2���4��
��(�|��5���L��z��pWlR��r�ɤZ����P��"L�1��c�1�K���֣�hFdLZ<!Z�\:�Q�SS����eĭ�1U�!��G����&�j�ǡ��~�"�A�&l�
�_�F�"��ÒT
��!6���@����ф;S�|GE"�$���k�:����J����s�A��v%z�,y%df�1O"x�c*Y��7�M+ydbs�紜ɭwN_%����v���'��k>	r�n��h(��	Ԃ{[�Du�j��
��m0�N�b���xa��6/�ٞЄ\�w�Lw�ͽS6,vG�]��x\�]
�xq�'��2�dH�˭�oZ5���˶8�A1b`�H �~(/�#�9e ����t�5�ѫED�lRs^����Rt�qOWa<}��߼C��9͂ �u�#�����M���>������e��}��c��މ��UbN��Z�wS%�#A�OpmD?���q*��3��!֒�y��[ B
�)-ǘ�I�J��;�Dک��b��*[L5�9��A����Fq��);���8�rB2CXbu<�Ng�(6���U�87be�K+�,�P~ypF���>4�nW��/l�.��Xs(�H5�o��(���*D闎R|�U>�B��&��4��U� �a/GE�Z��}��"�~�s��Fq+�6�A���Jƀ&~x(1&P<�����ˡg�����bh��eW��&��Pg>��
����[j_�u`�0Z\}s�d�Y�t x���O�Y���u�^]2��(/�3�J�D�eNg��A������f�fW�����N)�C��m����#�0�%��3�z�[�˛��j��fBZ��f
�҅T0uaA�vD��z��4�t��R���O�|��1���H�����MƄ�:�Y�Pr�f.Ō�������%<$#/�g�<�R�\��!=���U�ɴor���Ɓ����J��g=;M	��QD���|�AI}�Mx��T <]�f+M�|i���V�~��3��;�^�o�j��ɩ�<�s�PA�O!W����I�F��G�\S���,ِ���*�����]��9�ީ�;�}2�G1J'�b�����_��j��ְ �C>ܰp�@w��E�l[�,���2�%��H����G1j+��>H��O_���@����{`!:��%��nL��Ñ��D��(�а��!�qjP�LA��-����s-��IC�9 d���^qPv�w�@RF��3)���$J�&�E�oD�'�A�?$D�(7��~��a�!��a})�G�X@�;�7`jA�PթY@=��C�K<u�I$�	� <�R�_t�L�Z�/��PVzc�L�G*��eҖ�l�u��������L�)�/��C�s�[�Gq��G?J�x�uO��^i�ؠ?c�.e�i'��Δ���kn�NgO	�(S��H h�^^��e��wͷSbI2�����p��q��r{rcD��Z�x1��y�͹Q�o��J$�XGA��whB�6�6[A���y� 2�L�xɷ%�����18y���g)�D��3��A	��{i}Hf�=Ͽߤ��{ںWJYz��R�l���X�&.������}e��moU���^'F��p�'<�<���F@}G�w٤�������Q���/�h�FM
GcpM�P�76��κf�+r�ʂ�fL5�Wr��aj]�R�#kMXwW<���Ա��:��{�;IE�_O�ې�6@5M]+i4n����a�-+���2;E�u<0�S���rej�2!���(�H1��g{W�F� ��!H|��)�c��|���0r�6`�-!Æ���\:3���EFG�B:Y�&�ȷa�1c�*�} ��c�fB$8��Y�]��׎ⅷ�ꊑ�hJl"U"���~��"��)��������j�:���H�,���y��g"~�# ����wVǥ�z~i)�Ɓ�[��J�gٍ��!\gO�.tA��<��*�^�Aw�Q�'��}m#q�mO����)Na���d���^$`�%��j�h؄t�}�����n=ҝh�1c�w�6��./#�6sP����1���^�t��O|� X�y��G j�-��G:)8r����YL+�Z��tm�!-�:$��$\�IC��{�?��X�,���]�]�`ECFH��B�����(X��)��<��2��m:V?��s�O�w$�Z� b�� x�-p��M^�k��-��<�ܒ: ���-L�a��w�4K�Ԡ�y*»�a�g�Pk��0g��sT,��0��Gd_�}�Y0�����=�����[n����b����v���ˢdh��rO?�q����������b>T���@�r˅@5�C2�}z9�1���촸e�!B�Б��s��+��bh$u|�;bDz�(��Z�GWq3�F8XS�z8 6v�V�op�?��|�j+�WPl��c�}�!�91|��n�z�]�g����X�U�%�3����xz�G� ��
yT_��zTI�uz������U8e����/%��� Y��������jw�+?[lj�٨zh���y�JiPE�d����VA�N���b�n��Ι���0��=�|�/�#֙�T(���^����*"�8'ڑ����W��m���1�\X0zL �4��Y��C�BWX�(5H�-h�B�m<�Ύ�s���2�q!�HQ��h�:D�Z��i�ʔ����¸��0�����J���=�=���3
���������D�~�`R�W9��o�L���!Fr;C(�t	@:|D���`��$ �ň��K��jO�0�VH�CMG��_ϴ"��>YA���1�cy�1 ;"��!�N������O[�&�z�y���q-�)��<f���'��=��7, ��Z��K�CC���@[O��()C���6��.c_���vW�/o�yx_�,��?6���%.��g�:���9�e�)���Uekw'q�/宑Xe�+�T��*�,�x�!����O�I,��K@��
�?m������1�W�p�:�Lä����\����6�ҳ�j�V�|#m?]�o(�X����w�n��0ڳ��B�&��c��Lt��F���%i���EAi8��A�����U:�n�TqQ[{�9�Xk	��pD�C9���>J��n��� w{���fJ���rOҲ��լUW7���	A�Q�i��>R�_���P��CG���R�xt���8�X^W�cմAZ�U>��:x�otJh�A`��[�~��LA������
��0�7�jrW��bz��e��m*"�i�ZeMtK��͹t��_������D���`�Э����|۫99oM�mm���T;s"U@�Z)�頷�AcQ��!ɩ<�ۯM�a@jm�G&x�/��湢��!N��w�ёv^\=K"\�$��A�?P�n�V�;��@l��YL�l�K�xa���k��>n�2���
S�ܪh�~	�Mπ̙
�q�R�q?٫�t5�Pא�F������r��!�������ׇ?6@~(��։�t�:�y��I���X1�'�V���������n�^��
%��h#ŀ���P���U�8��U_cû�/68 G�|�a�?'��L��"�p�'7[Wq8������GI�9I�(홮��uL��2�nV��eom	�����Vp�Np'[�+j{�?S���t�5�
)T�m��*dyts�|���`�i?'����+��g��D��>HH�2�;�R7�Qg(_e=�2��°���LI�2:-?�|���?�2��+u�6�L��PFnR�y��P��}4�݅%^���v��[>�~X�h5�V����2�"|�`���>�C���¬��/����`<e��m[�V�L�*��y����Ӛ;�\�R?�@�Q�AJu�������4�w���R������_�DG�h��f�U�\���l����ꨄ�fkE:�#��X��:7����:�CnCx�OFIH�9%� 9���O�(�KL�/���bxH�EˇHu%�G�C� }�o+d���0�ƺ)QR@ᑏ�G�1��z��ܦ$�_�Q[6�����&����Тo��Y(�!G�Ŗ���XE�G���:�ڲw"EaWqU���F�al�׊*�8��#@�u��B'.��VO��ar.����iB;>y�r��jGmQ���LXyi�
cb M:��ܣ�C �.yO�K'�q�.�u{l3ZFA�ͣ��G���W��iG]�Jta��~>y��짔Z�|�0b}�����q%\��h��eB��1�RuQR\u��D�,ϙNo�n(���!FAI�ܮ�l���3_;��>巽14آe�
��h�0�ĔehA���$�g�kAҹޝ�脩���l��*\���L�쥪CM�#��̪d��RO�"�zO,��JT��U^e���vr���p�c��ɲG��E�����iK#˾���ٕ��@����!Dq��y�N 7���U�cg���҉[j�����P��T�d`�I�&_�E��l��s[{���8����� �c��!k�em+zϙ�<���ƯX��ɪ}�O�x�&��3޸p0��|�Z=-~$ѭ� F~R�F��n�b�VTɯ�F�<U��+�b�F�G���W%6U�k��-���*�{��ک~�q`N����f� ɰ	�Ǘ�W���vT���.�Xn����'*�B%<��sXHh�<��.-����mv� �l�'&�c)e5K��/��I8���,ܕrf@f��	y��a!��JX8i]�M�� �i�Mk=��_��Cf�V+������O*k��b�[�j�e����G4>���j��a����&�/lw]�ד����,��.��NyC�J8O'���wvM�s�F9�״�󻡳��}��:��!�_'�6�B>�c�ƶU�e}k����;��[K^(ٕ�|�1����ە|�B+]��d0T�`�U��]	��$.�Hd*��7�G"�D�ƪ�cƗ9��/�ج�Aڽ\��}���F�Y����kC6�q$�����gJnsk�O��� .���8�6I����ڂY��P ��%������ =]�#=*J����߃]z�o�?��������Iѝ��c�5�tq���V���ʻ��p�C�Ho5�ؑ~�M@���>53�-`.�-௎FK�]/V5���Q!mY]�uN���x�@�9- W5��_�@�K�����{�� lZ�9��P�2It-%خ].Z%�ǳ�B�A� ׊��7��ރ3l��=Q�|�� 'w?��#�C@�϶��Tk���Qi�p����/0�6�2LZ�~ѱY�
mCp��t�R4��wo�ki����4).4ۺD���&#6��mP�|�s5#m)�#28�p�����ƫC�3	z��Y<7�@4�R*��u���!f��B֒���aH�uPNE�[�).���i0�B9��m�!R�C���I�y�qFkB�}���#n�<a��~�`� n��;������Ij��%�5Z�0��	��t�"��ӳ��cmڛ�Y���O�k6ez@�/)[
�{��:��Y����B�wABX�
/J��_U���S��XaS��ռ��i|�P9�
��YdA���w�8���5T<聹lj9%0��B�
<R����T�7�HU
���qR���<������l%oN}����	,�a���!���j\�9�}k���ѣ@K��k �c�U%�̢��L�~^ F��%�����9/ĉ�k���l�`Q9��b�Ϭ�IXx�f�|[P�JW�S�ڊ�Նq#�Us�<��]���4����9���q��b�+�	��^����{�@?SD�-8,T ԛ�֟0���XOi�Ɨ��v��B���^���u����y'��>�o���F�4���j"͐���t	���E��҈<�����R�U׷9�Ym�� �"_2!$Fqkr��| 4�,8�r�^����E@E&�5Ҩ�g�o�?yq��U���&9F��El����v��Z佱wAo-\��#���Po��l�/(˖W�Z �	v*C���2���z�ܣ,���:7���G������#bT�PS��Z��rP	Jlö�ЌM@51=�\0v��`�)$�E��T��S��h_��N)j��BJ�3�����J	��u�$;*K�X!�#��wh��k�)�+o�Q�ٮ�Q�u��`���*�Mӽ�y�BYl�D��M��6�g��U*�t��	_L�Hk��~A�{<�X�WO��fY���x���G�7<���
�D��CMEt��FƫAL�׌�� �n&�~�T3�.�@q]�rwK���\��㰿װ���1�j��Rn�J��O�C�\�*�Vߪ�� AEKY�{��U��� qLF,��\�(��ݰ�'�%P�Ѩ]��/&X-��<��e�@ܢ�=k?EH�v3��nS�ѠLf�i_�46�^l�9�5ހ� ����m>Mn�{H/3���8�h p��|����y���U�4�[}
���j��� �������2#�<]����t��|X7���~,.�|^����`����9�=_�ww�B��M�wx��5��7�O��h�v����bh�r�]^�� b
���������E����#7�6�ǡJ�n�<w)?)��|k�Xw�X���xS��$n�V��{\��L���x�9ܫs1W3��(5�X�w�w����ʢcPMU���x�)��~�Z��7?>�L�5��e��Z�׶Њ��b!I��+cw�]��`�x��t��	F�C��$��aP��+��+��'R�n�Z����0����hq�RŜ�s5��N�����`J���}8/Mh�%%y?�k�ó���-!��I�EL-��7� x�h�~#��(s����S�J�xy��ː�]1xծ-\o�
��
�5�H?��]ɭ��f�}�}�hxe���L�v#o����p&`��Z/g�T��s���h^���?���K<�c�$Z��TRlk.!��򕓚V_;��z�x��,����5��mq��/;ӆ"�d��m��4��-�$�H�]Ru�!��̰B{49/��i �%O޴3"מO34���7(�L	�'ױ��	�l������?:���u}?3C��U�ؤ��	4(*`ÅR�K�2Ҿ�Wy;���0�L>�X�]/��]F���������Ŀ$�� %i0����L�V��:#�����%KyF)�׏��=�h0��'�K�h)��2��ѵg�G'�;Ծ�A�2�#$u,�iP5�U���g���Ίv�̭�l�!���)X��Q�$� ز��Q�NR3t�!��-\u��`	#*$�(�[�rqY��_-���m���oKS�%�L�W�6��"��z�Q�ޔ[��n�؅V�+dn �M"�h�X�|%`����6[0�@Ϥ�\����	ϛ��u��g��֞Hً�%��N)����X�x��A����5X��������Ϲ��eg��uG�kD��G�@OY=��1[�L9��h��\Q�߻��B��?��qz�m
 �:��ל]����	���ҷ��.w`:�'�L�>_y��x�#3�Q�9�9���0$�� 5ُ,�� �FP��<����ĜSw�G�����X�1������ ���� ��!\ v_o�㬗��	�c���?R@vo~{4aQF !#���m�y ��V���"e���a��K���$�o�Q��0�����|�5��H��<�=M��l;v��g�Q|"X����G���^�@ ��9i*-���|�D���᤾b7k@9��r�Nd�����=z̺߮VG`KX�C���d�rѪn��JTG�2�w��_���
��Z������nؠ�q����Yt�����W6Y�ʠR7vK���'���46s4����v����߇����J�j-%���(� �n��ǶZ� a����W��'ИC�Q�3K2$(�:����^�ٳ�u��X�7&�`���.k9|:}j�i�����M�ؖ�c��O.��O3a�>��}��B�������f��$�CG԰���qX��E��d1�5�� ���zaQ���8�6\�V"M��=��EOe�Wo���u2���"��E����,@��D��t&�1"��S�wK�p��E���eN��u:���Li�T��d1,<�	R�4I�|�4;#���r{A�)j�Ad�;��Wl[�3�	������$�x��}���*c����˼��Hdul�s�"��j$1�׼��C����ؽ��I����U{1���.�J���j5W�(��$8�Lb
��/���`v�[Y	��d�����&Jл��824���n��:Ӫ��Hn���BЌ�1;��`�r��h�]E�A<��ԧ����(��fأW_?Z���)7�T(b���c@i���6��Ud9vX=�g�����hs#��i���vB"��`MzY�$�"��_�p�@M0�boV/n�gn���oG"��FS��I�"(���F�U��_##t54�nӨ����9�79��a�a|�hh���T�3N�rS1���?���nj�����M|1S�?�&�Lj�$�F2�+���|0R<�Q`���8©���G�����`E@���/K3eA�����%�����%P�S��ϛ3XLE){H0�3J���LQI�
6۷_�<T�?���P)RKDؙCb�*(��Ő�̿�44|2��	ջ�,�w�z�Ag<=b�cx�V�̵���l��h���osk��
��	�e�����\@��^��O{$���`9�w�!�BŪ�I���st��R"m��V�+�&d@��]�I�p5RT���^�]���~�8$�,zT+ZqF�	_�d�[Z�r	�L3�ъYS��P-����C*�ܧI-���:������`���E��]I$})b)���"��#�l"���b8DogE�эq��V-9g�~��V
�;|c��3��ԙ9��!s}�Wp��l.я�ϲ!]�t�	h�9�dᤶ��`V�QU��;�9���m��a;��F�A�$\H|d��5��n�0d�L����)e(ͽ!4�t|.�����|�
Q�{;��Y=�{AsY���]�[���x����mf�����b\�{+ɋ����AF��l�'�`�[#��+�g����&c**��aa}�_4~�B�c�;ꅩ�[N!o9?AWfs=�-{����i�A+DO8��V1��:�g�[j���KNU�&
6��+��7�a�f��U~ފ�b�-�6�i�T�W�5B����U&�yT���_{q����@�e���om�0�9 ��l�e��+�m���5��̴97y�Q�"�g�Z��a׋w2�n���ݬ�P�4ZN�������⠊�-A��^�*�m���5��[���l����m]�t���6lה�^j�-4d�@�t|®\�c����	� ����~G�}���T�Fceڰ_4�e��)+�^!�~'�k��Ƞyw��\�%���&��&��4:�������<H����P}�t�ҁ�$O��u{��L?�����G���Sb�a��p�_�4���l�*f�I["��H�XGߤ�TƳ����QL� �^��U$��YJaĭ�7o2+�/�9�s?��N\��(!T��H _o��䗈�JiQ�@:��<ȶ<�d��J��
���Q3鬥�s'��a9��<���<����x����k�k>F���7��ݬ�V9�O�SD���Б1��	�ƞ���)V`Sj-��e0�J_S̀���{`Cw��W�@���p@e�t/=�5����I�1�ZX�a��X���p6�Is=�8����^����Uc̟�eq$$l��x�o�XX�z����i:R��.�e%Pt?��s���:���r�����B���ғ՚��+��"JO\O-O�±��*�D�ld�`�i+��a�4gw�>�6Xp���F�(!�:�=j�� )7�Гӝ����:���媷?P+z�KI��p~
��Z�L�i0*�26���ny�e6o���ߒ�,�5r�-�_��n��`l%1�>"��zXp\PNc�&#X�8&�u˦b	p��@�����D�pP=��M�V�>6�_`�y��:�Ŏꐯ9�v��Vl՞�d鷑�\�ؠ27�U�m�@�o��G�7��'Д��D��W��}�
��X�-k���#t�Xz˹#���Vc����#-g�SI�ώ	��M�&Ń����B��r��r�f^080��<I����7V��"��эF5��
�n����_{ϛ�*O��@=2�[����_9.����.�y�@6нm�Z����|ȥ�%2h��6v�I�3�3F����h7��͞B,�Okp�q��n���V[�(��	K'`?�E��-`�y�=���g_j���p]�-ϑd����,���"��E 	%�pƠ(8�rn:?{����?P8��G&oe��U�6VU<f��S{��wM�����:�^��z�N�q�ڛ���l�W`3�X�p����.�>7�Oz|گQ��.) ��ˠ�9�vqSە���4 ��S�J��� 5z?��FAy/.Q�<�������#��ߘ�-�!"�g��>��+�Lz�;�m`�\맮�xLm��PyhΤ0�q^���P�;nP}j]M>9/̓��;�	��б�m:�����
d��;��2�x���k�+����[d|�	pxn�i�`��$��Ijf��P�D>�6��E��󔕼��q{�v�ߵ�UW����y&�
��T�~�>�Vq�&����CF>l�a�d|�GJfی�:C���W�F���v��.��n/����QzcBUz�~�Bg��YF�{��O%�_j�<o7���s�
E'ઃ�C����B�ܮ[��^��vh����Xh�:jnXqQ�D�%|{_�`{�G���������8Pk���B�;5H#&4��|�3�A� y�BW���q���K��U��Ȕ���./�E|�WDQ��CznZv��E$�.�ub ���ܹ��g�5p��~WD��1�# �I\XS����Y�����0Jh���(!Nn�*>�r5AQ�n�����ZȂ(�hp��Ҳ��(5������c"p��i+p7&���z�\#��4c�5z�����m�I�
h1�W���ko#,"a���1�I���N5���qx.ؤ�� �`�j8����:�7��՗��Q��Q�m0�}OyHQ�S�9��@m{����
�I�!��o�=�H���6:-�:�
X������;{D(�s�ίǒO�s]5}�͘�ᇖ�(�'��_R/>ސ�Դ��6*��$�C��!	�κx��U�|2T�ѥ�M�62��X�;���ciX�<N}�Jve/q<㱤{:g�x���u��cV|bl5\v������eA0K���fw F)�]��6ͮ�o4���԰�F$�\(95�0��4�~�We��ȅi�rf��b��|m��/�%yj���^�.��|�?	�:^�������N��%�b���x́Y�i宽3�@���Ĕ�W����l���4a��G;ћ�Q"�v��ȷӬ-�?�x�ʢ�ck���:�y��C#�X�<��wE�?�"�]� ��������L!���g;*�b��\�b���e�a,���&n7�隴a�++1�j�? @T)�W�t� �#::WV�6�rl����y6�K����K.�	��r�"MԾ����㡂2B�O|�ݐ������F���k������:t�.�ɷl����C8e�#/D�������3�/�N0Dd1���,& �W�M�����V�����((�'�(jm�L���/�oY;���9_��<���x}��>]�nҷ��fw5��t;ݪ��.[-3���M$$3M�R��܎�nt�\/)�K���s�3��A�*�����p�k�F��M��/�����Yc��f�4�����E�wH�ՒVD����q���|��m�:i�Yo{Q�3 �4�<�೸%�bY}`����z�i}\yj��3b96���4J�u��p�l��U�	���J��h�#WT_�#]�,�c �B���%شڢ��%��C�]OR9m��7���j� ��"�(��s�]�f�1�޲m�z��J �V=�-aG��X�O-_��o���y�YA�u܊���&�C��>'����1@�b!����)�\3�4�p�C/R �����ں^�&�:s8�_��0�3��M�N�,�����[�״��.�N-��Zs>3�'#��P�f�f�]
���}�&���$�[��tD޲�-���S�?Ѽ1Az��*��j. Żє�j6�^T���O]+F�Z%�4>��|qAֹT��#�5�0b]2��J�}�HF��,�VTC�5I��C���d����[���u�P�\��8��W�彁)��@+V|-M�z@E��^5[�������������O�8^�s�a:"��Ϥ|��g�9U��(H����`#1,��ʪT�v��"N��M9����M�6��m�m/&�	Ne��[8��)��"p㵮T��?v�3�݆�w%V���pJЅth�b�<1Msz-��!����*;V�� E0rIZ�$�+BA6��u����k�+b����v������!o]�(i,E��KR�M�:P1���+L�ʷ�9�m�EL{���u�<���s�,Qq� l�R�[���tT�����n���\lY���}1�8�fdx-���:�p�mdw���Eӄ���3uc���q��w��wJp`�!���	�,w�Z�;�d����ݘM��ۻ��f�d���y�!'����tZ��I�b�{��7��og���� 1���.�&�'n�O"�Km|�џ��W���0?��.�������n��2�iܕ��U%
�<�"���nNw�������H�!��ϧd��v$(����)ś-G�v�#JyHC��լb�ܔk�,e��P�K�O��g�1 <�=1��7�[��D���a�oT�A�/Df�S}�㜋a+]���_�VǚU�SY�d��J�?��A#��8M�>�\P����O0կ\�s��Yj������1M�������,���sf*7Mt�L�%9�e�1�U^�r=/0X"	�A|7f��_&-�|�@V
m��_k�vB�vE����$�'S�_`Gs��EPŎ2E`4R����}�����c���O�OG�	W�~�����0�Ig(��7�u����C���#��g�l��2��NlAR?Gn�r)5���Y�6�Jϊ�`Z}|[9��#�t��غ|�)8�g�����b���g�J>�Ŕ��� ��Z<�O=�����K��h�5�{'��ڠ�2�Z�t�>3���6����f����1��;��J�˄��9B`���j�`u��9#G�q�K �E�XT���Y�I�� �B�Vwf�.��,3xϖS!��H��2@����{F?v7l ����}��a�?�(X�,j!$�n\V�8��4
�*�F +P� ���b-vQ��ȷgK$Y.Rb�:�J��IN�N]ڕ����x� �L���ʡ8��c�i���^1�k���-��X��@���j��/��M}��)R������ԇ�ce��t'J�y��X�@�o��T��`�K�ɍ�lF�2I	���]5/st/��P�k9etPPѿ��"o�[��`f��>.z[w��r�2%7��,�w�h�
FD����O!�t���Z�ӓ����M��U��ԝ��vx�zWC;��`�`��	PM78�M���@���r��?1�d�|�Y1��0bo�2��}GEީ�B��j�<yL�L���	@H��O��VtΔ�a�"�E�D!�g��239�<oBr���$x��*M�X�sا�ʿ�I�[4	�~Cd�a	p��g<�qB4�w���� ��'�����b���x�=�tY`=�l4�	��ì-D��L
:��Ǧ����
<�z����[S���Suٍ�6�����~�����;wJF�#o������]5�ɨ��i ��I�]���?1-.��[��WŻ9_��i�6@I�����e��?�ktL����2�3׉F,F��J�'��e12r�?����*����êr=�JeYA��y��T�ZӭC4�����`U1�9���_Ì�ɺ�J��(�%��Y�h���L�׉V#����Ԉl�q^��X5
lC�m��¬�����ه�j��}��4'��['��Z`�����[���u�W�o����� ��ۯoZ��""�Ɍo�%�G�#{�:� �|#J��/���N�w�P>�hs��#S;ҹմ��Y�M���ϔ�����o�؍�sc!HH�T��f�u�\�!�gg+Y�z��T�~��!�tE����T�9�(�4��|�N��yqd�~lL�#"���D����!]ۿ�& �|����A���'��F���t�.��n"D���R�m?��1f��t�9�y@7���9��R���Jkq���ƅ`�<CP�V=tٗ�|�J>z`��]�;���?!d�bx�<9�{�33�4��?���ܞ?n���P[F|z�$}S8�W�j��s��������iP	? 
�U�u�6(j6�C��(ZKs9�A�qf\C��5�����[)�7��1�Af��uB��+��Bz�7���r�d�������CG-*��-��(��G��ž���|��Y ��h��� \Β��m�5�>ܜ�Q�@�9^tćHO(*c���IO �/���fV�f��T�M`�ʘ�u8��<A���9��\e�0xvnXé �YέVl���
�n��C��I4�z0�C�F���n=¨uD'7/y\�X�M���N��O
��b�W�Hy4i&�'sm	Ѐ���z�*��9�c6b8�B��X�w^�����!�^aZ5�z�˔�~췏*�X�م􌖞&PS���55��'mtZ��_m�pw�퐩��U7V컊W\~�|�Z;�����>�e�� d~|��pڽ>�;Q��t
�w:kTa��I>��v1�ճ��z�DA�1v@���E�?-���8?:���eW�J����^|rX; p`YN��Ԑ��E�BVY,4����<��Ya��	�|�aB}��h�u�|�&%f5C���Ԑ��������S���w_�CUy)O��8h���J$xR�O�hD�g38�����m���o��Eb~�'(cx:�v_�ײMc�!���:`�u���_��.K(q�H18�ۣ�����6���@J�R�Ŋ��iZ��b��\sm�����@��U	ʦ0�.2hZJ#�	-��t�;��C�~Q,?ЃY�x��"�R�.
)@�:"ĥEe1q}��o�1�e���N�4���7fj5�ԝW�
c�ϩm/��;��Dy���~m���ė�/���<�
^��3V�'Zn��kّ�;�mg�nAt"�'u2n�	�љ��5�6�B����V���A�B}�=^9``!��P�)��k5��Q\�Z��[�@ȉ�`+*`�3?G��%d�d`^�o"L���FXRD�i
��7C��'��G�=���s��&�&������jG�9��)b+߫�r��j��O��i�gC!�D�1�_R�by�V��dP''
t:���3�ƭ�#�#\���V����E7Nܐ���ud4{̆qc�݅=��A� �h�X�A�:$Hn(֫ ҩ���l~�td?�ހ8�j~ҳ�ʀZi������h>{礨10�Й�1�4���������\��el�
P���tq���^�/���3 P�Y�����ÅEWA���t"��҆?��-�>JJݹ���r�����k??��.tB���<GO�
զ�5�?�p	kك�������
"5ql���q���L���ֹ��Q'S�V1m�������NS�KMp5�:kSy�7A7�Q�#�(�՗�W?$	u2t4XvFwJ���Y�NP�D�V@T$Aq/
�J�h��3�8�7��zmA�9�f�0�lo������<y�+����;/��ӷ�n$ic�V�$�X��W�B@��`*����� �6��&��)��Ԇ��ë"�.�<nK~B.��$�4��7�F��Gah���T���\��E��hSM����J���!լ7�}���zK�1��:M�yK�m�L�q�2+Nt��3�j�w@��*��}K�m��_Ȟ1�F����M��Ԛ6��C��yhk����E��\�86�\�n��o穓V�kT����葕-R�[�! �^C]�ͦ39��=%���;M��}4l����E(�>��2�n��	H�����{J���Xx&'�F���ܞ����)7L�3>L�}��g���߹C�|G-�Q�X�5=�E�����y��b@�pD<gN��[7[��Q�+��`�n��5�p�*"�ZM���\�h
�hA�ΒaM6�%���ޞ���-N�:�B�U#�0�4�-��x��H¢���/�:���Т�}l^K�{HU�$L����,�+zw��+��|���-�K��y �!P:������+����f|TdH=B� �,� s����Z0���䦮��;��Kΐ��|�
�����E�-ޣ�nI�:<�ӄevY�b�m�l�+��j�%���\�F+�ʩ��J.e1Jo�������E��"xv^*M�>�R�c��Y���䳯�&'�� "�O���:Аۋ@W��(,�sX�x�\{�}��ra��L����n"�Wf�����t&��4�y���O�K�/?s�x�F_B�=�L�o]{s�r7�K=p����j���}ۏ�$
Ăj�xaF@ʚ��nJ7g���nAU�k� ���q��<�r ݏ�pK��p�䪶�$����e���$0�-�=�6�!H��0Y�3���������Lzgj2]��_��v?�H�4F?Sab��Q��8�h������O�#��ވ" L֍�S��/3���U��8�f$��'/����Eםv��8`����0E�<+�88M|}`���
d�����3�v��I����T*<Ʒ��D���x���TY䌨��u3�T����V��'vpr%�iЃ��1uo�fcr;�۞~�|��gb|��p�s������U�r�����e3��H�k���k���hZy`-����N��%7���G��{�2����&�iSIʝ�$�]�7�5� ?$�\Ѧ����t\qe2�	�N�F�b�}�>Y��D�X}��E��cߙ���y�NGה��6�F�w	Y>����w��5�-QN��$fK���^Q�D��1���ۓݴ�N�� �Ű{�KiȰd��؟�	�o�`B��Y��];���T�/ԇ⚉�����ͮr!�f_"h��b�W����ws�=L'���{������u0�Ć|� 	+�I
�\��b��>�o���F�j2�%A���]��q4:0Z�@�?�d��J��1uVy�q�$6��p�M��#��v���6Ůx �b_�;�7��LQD��Gq���?@�
��g��0����Ցl��I½����������Φ��'.ǛA�"t	��I���³��`�V*&\��n����A�y�~��NhR�È�bŭyX�ց���/��h�^𪧖�/ݿ]A�FE�C-&�RYF�@�����IR�&�S�C���hC��r?�y��� h�RUNv���o6?zz��Hz�z�<+M�ęM�E����DVO6�Zd�r#G'�0��vvG[��Q��L̺��\	t�T�sC�s:�RQ�D��T|󣾮���QW�a3e�O�i�ZW�	GՖ�z� ��By����?TFˊ��*N�o>�vs�)^��lQ����?	��s39�a��&���6s����0G�^�_t�6�̛	�X�F^���(»VsN�!�����f�vtj"�\&�v��}�z��`9a� 汬��~h;�6av����[�?./Cǭ��?�����kA�A�?В�4�j.�CI���ke��;v�x�ˉ�g�� 1�GZ��#��Vq�/V��JY�ؕ9���GA��
�
﵀������vɻH�NV�zް�$_5�.>�c�s�E��eynP���_���j� G�7�rc8�!���^�Y{ɶr	�(�6�e�[�B�^$�[���
� iS�0�i����iK�k
y��2��������m$Y�<�,%o�#��
)=TB÷�,'78�i�T�>HJ��y�T�����:�'̼�e��E�"�k�|�#�%CD���_�0���m@J��S0���u��:�;\+=S�3o�84
��?w
�����L�]���'R�z���yr��C����B��!�J�|8n���;���?��9�������D�D���:q��.�X�dic�"�n*G(R���#[T(f�� H��4~����2��Q���#��m�X}c)V��>�=����n��"�V7X?�ˎ�����>W�@S	�T�M"0F�R]�J��0r�r:Q�����3���MK*��t��:=��i�.H_�-6]QYuFC�H.���Q���P"�n��T�w٢� ui�`[���[�Ԣ�v�'y�+:l7l6�X���0�+�����ZH-��	���K5?#��/�*�z��3C�sq�m���ln-W �G�p�B���3�����xu7�-w�l,-�m�R��oY���Bu}8O�kHx��(7�&���
�2*D�����c&��{v����m�81�v���r���ϴM��d�H��%:�BCE{���Q��"7n�A����m"I���c�Þ�*�TA@��l�>�vT͞H(�._�' x�����#x���ghGO�'��G��䌏0/���8?���HP�r�;�R�8L�#-�5����)��c|b�?dr�LR��3C2�m�]Z�ڟm5�ڥ��Y���kj?$U���cz����N�Đk��h�=N�6i���z�IdP��YVMxZ!ods�7k� ���c������w�Z_��&24.���C�uE��.a�P�/u��[����յ���� ��Aj\'f�+�SC�cv�2��N>�|'���d@�K=��0��8n/گG��q�HQ:����4!��2��Jv�*�w�Ǳ�*��F��E��<�x/�.�}s��NF-�#!�ꟴ���)�����F�{�q8bN���H�K��@������?��\@\jU�]�Y졳�ظ�����&��#SK	�:�U�7<��nu��n�^	�0��_n�{B͜+4��b�.<��I�o0����LL�����W�B��9��Y���<�r�v�	�ԡf�Sa]�op&�,҆ĩ�{%N֫h�}$\h�2�FB��=�PF֋`��u�^jpK:>�����L��bX#�J(���I���K�C�y�6�5�/T��ϣf����n`�=�5�m�b ��/�X�a�E_f
cV��I_��:�4}� ����E<x�']��>wQ����`Oy���8s:!�z�:���d��\��D	7��a���I�=|�&�\ƌ�J9`>rH�^��I�n
�ngk�}aG6��1�o��8��l;�|�����y���<Q���fX��G@W��r�]�l�.��`��rU	�.I��}��<��B��1S�h�Gep�'�C�7.T�F�
�N�5 `��Q��I�HJ�K�EL�:�[T ��6]jk�3k*J:D�,�� bh�n��e
4��{]��W8�0��ۭM�X��(Y6~{�*�`e� �-�KYL�ی��ФW^C���G�4��8�E6���j��G�yX�u�Jgu�:][v���;�w�����w��s�8S���۾�5�_ד h��tl}U�v59:n�����9�fUٮ�e-D�GZ�D?z�94fF�@X^<��*w��+��p7������Ls7"p�:����b�y_��-p��g���v���-\��$�����\���CȎ�y��i8Շ�m��^c�vյ�l�-h��e"E�E(�<����m�k�x3���3YR/N�7��'~����3��tы%Z0�?�c�����6�?�;]��C	/D��q�wn�ۛ�%ޱ&�j"��
���I*�z�U�����\4Q.������#�Em��xc�Kt��I<����TM�Z}�#���oO�)������0�O�P�u�pYȭ�F�3q�4���&�<c�ҙ:�G���>;���P ��Z0;@5F	��^*
��J_��|�K��f/Y�������p,�%kT`t=�t��]�t�2��>7�o� ՜
� Dkb:1�y����0����f�_�	I�V�-7R�y7)��-�@�[sK|�ѱ\Ȕȍw��3��������ěR.�V�{�0B��4,�WP$
��M��]?w�3徖�Ě�7k�e�|�Į	����G�-�R|�Q�%m �.7s�\�8�9�.��ce�S�I-�:�����w�9�M��;^�Ա���I��0������l�fY���#��CH�V5�eB�ī��u=E����.����9-3FV���z"P�
�P3yzR1�2t�!2D5��"4M2x4����|B��h��	ds8jt���ݜ���(�g�k<���)⍒�F�;��$o���8S�G��7\�
���� P$6w;{6���I�絴<�}�u~�V��}��Β˳�I4���ԭחEbf�j��!o����#���Nu�V���}KՂ9��u�PJ�8R��V=�~B�6A�y�_7�ԹU��"��z�F��a?��A;���4�p0�֐L.Xw0Uא���M�T�nYcbo���A�qZwc�vӕ�ok�h.�Q"3�57�]��_3�cr��I��C\��se����>�����W���:��9~�D�����*~��I0aL,r�Nwߋn���'}�N�]b� B�	���	1b�s+C��2�H�Ůo�ӵ݀��a�/�t��[p�Yr�pN�%�^Wó4X U:WX��j��g���`������V�i#�x,�c���25g8O.���%�J������㨳�:�M��0/�FkN�Ry �E��.� IZR��Z��wt�W#([�}�^G{Bj�I�����t��������LKJ����:�Vo�4<.1���� =id�B���V��K�<y�#-'�=��h(�а�2p|q`���4.���Ka6�<@T�BOn�on��[�t1F�N�(���&��A�.T/Ɩ��$k�J�Ƀ����1!�he�������IS��B�s�}�Ճ�w���m�5�'=�&�u�X���N�h�n+ø���4��B>����il4������v�F��M�B'9H�O�L�"[ � {���r�VC���pi�=���,��kQ�^��Ru$cH$��ZdnAE��;6N���'c?�(7Y$�p���C�!N�:K�����)J �6������ULz6J�a[�����0���.��e'�<Q�9K���^�5l���@@+���:�=MU�e�^�q5�R ��)�;7D�Gmn�"�!�#n�0���۰��>k�0��v�BĶż�[F��],K�_�D�����4������;(�O��p���[Or��z�4 	\��پhb�wm���1K�BR`��sEZ�D�f���
�/��!'��M��K�n:L~Q���x��.�ž�z�RS�f.<�N�2Ke6�T���z�y���rGC���&�iX�F�����挊qP<q�C�4*�	�CA��t�\^��P��GJ#��n���	���S��tl^��/1IB.����v<� 4u�q#�������#f�ٓ�OČP�,JV�>j�,�|�Jy�� ��X2L�G~8��z:�0��-�Oq�i#��GzH������v�ӯ�P����M�n�W8�8��?2U���5^,u��	�(��tUp�o��r��t����7J���K�l�B�Xu�OV�{P/��r�ϧ�U�)Hbc��?q��iޔu�əxF�Pa�F��t�{�2f�	�i�;���`���^Nu��qv��kZ	2ǋ6M���َU��I�Љ�L�-q�^{́E�ټ#��ێ=�6j�����6�5<+���yw6����ʊ�Ƭ�o5�q]y`ٞ�g�PJ�e�S�E�k����|�(P��H�J��D�H�t��m��*�N�ᓝϖ.^�b�̖%�J¥l�Ιg�M���-�D�D�u�[��'c�6���c]쯕'Ң�;��|/L�fX05�o�	@�vѺ�:��`\�ק�xR�d��.H�-ox��L��M�b� Q��/	0W�E	��crz��4{8�>S�ꆄ����_^��D��AV�W�b4�4z4���a�cM�m�PNI�q*uz��E_
h/�7B9tj!{���4?�vU��N	B��!uCi��m�c�7�g�7i�%�F8V[��j�ᬎ�n����bhX!�C���z���-4�=�\�A��);e�a��Æ���Lm	�#�pX$
dO�(�*7��J33�~����:�v�vRL�T~��ߙ����1:�0��nC�1<O#�5�H�Q	�f�P�_4������ ȼ��Zf��Q�	��S�NtH��[X)�p��W�[p�]���u�X�@����|���GR{r�u���/�^�� ں؁�@1ݮ���#ʪ �Pa�D6_W�K$�E�޷d��=GՁ�5փ:��h����Bv��S-#�w��9x߭5��]|*B����t���[�����L@�u��G&6U5ģ��OM���nV����*N��Ö��c�c�A�2O��}v�B��۲��6� �F����wZ��'�S@���1�������d��Jµ��g3U��oo*�Ja�ey�Q��H(��Ƴ,&r}��X倚�C�u>�fƦ����9�l'R58k��󂄇3���L�*�\8��`j�MBI\�I�q��O��O�׸s�Aܩ��:)+n<:�dQ(���fc%M���9�G�����o���
��n�S�(s��U����,�/�h�\�>�D��4B�l�t���C@����Y�UYf��]������[��w=�5�<Ș�vUQ�۲|)")��i����yk�03
��j��{�V}�D��l��nq��7o��fA5
.��y��"���53�kg��xMf��M�V�K�#���b ]44�ֹ��|x������:�ZC�8l58�5}��<��Mw wVw�t����`S !{��x(�o��ag�ᵴJ_��d�ӵ�2&��'�=R^�V����	��F'�6tH�AM�����Kyȷ@+�C��`0p�����/sqk��ebT�P)��95�L}I���0�Q�Z���i�׏���o:�q�D��Z��H��K��]��w8���n]y��7_�F�MV�<���� /S�S=��W��G�hцhi���nq�,흓*˧	]v��nώ���7Zy-}�a�ms&Q���������B��l�;t]�28!^���1���"s����]EI���Y�@�h �h��� �*e���ƍC�$`�W�P ��P�\0V�21]�	A������X�!�]3�����F�3�.�*�&�D@�K-gܴ%`+�_Lֲ��)������E���<񈭇<n��*<*f�
B2
��z��@��o��؞
�ُ�^_Ok������Uc��ض��4�%��'"��*0�Y=���M �3��M��oG�dBl4Z�q�SrQ��N����"�QB�rn��F�>U�&���W{�9k�Xl�I��SF�R�+�;М2K�!�ӯ7�6p~�^3۹��qgJ�B�y���q��HT��q��/Q�J��뗪�s���ğm�]`Ի-k"��F��AL������.Th�rL%��N�p��D�}��B}v�&cX����.M�8�|�T��9Pv��GT����sR$1-�F�[�I����Pp�����
͟���A�G�l�_����W�# 0��� _�d�Zb|
;h�_��	��[�����7&,���?xcң��a�A�|Z�j�(�s���Q	����2�)O-��B���s+m4�ё�Vm��\]V��^ԥp���:�Ň��������<���<>�q���`h@��/�yb=�}S��d/	
�Jt,��,\ISm��D�Xm��c^��X��I��k�����@[�&i6�L�Dw�� ���� t�3o�>�8�Q@mY�Wߵ#����x�	�u�߳�".y,�=~_J�����6��N��Mĺ.���:DT$�$:*#�c��	�:hS��À|Ezm��?5nF�Rv4��Q�����+u����xu���{1>l��i�6��[i�+��<F���\�۪Z�h��ߏ9�(ZG�����F���gU6	p9Yk�GQ��e�ĴW���8�J�i��k��w�j���M�'ڙ^C���S&� �\Ah���ý ��@�����,���T������M�A�T���p
����U�l��c�`�5�.iM�]�>T�����S~��/w�י�
�	YB�F�w��_��N����nX��l��X*���i!��7.�2���M��x��DHd��� �@B��i��	G&߸k�^���<�ۊ�1T�V��ڡػ2-Cu�И����%�ղo�q�e#�P�e�6s~�)Tǌ��B�*Y�<@�(u��.ʎ���0O�m� ��r�.Ȑ5:���Y�q���+��o��I�䠹�Ϥ�E�)����������fPrt,�ʗ��#�� ��i:�Dr;�w'���}~��Ĩ��HxU(�?�Z-\��Ұ<6�V�����v�F���
?��(賔Û��ʥ ����р����,qa��ǲ���C����~ی�U�8�u��7��W�-Ks;�8�_-fF�~�!�T��l���1;�$���_����O�����JBŪ���5e���UL�BwA�I�Vh=�L�od�֤T�1���B��T`G�q��xu�&5��ǫF�
�i�E\"��$�S>����2��#�'�N���z�ÃT�ܱ�!�`�t ئ4��u_������0O��E�(6��|R����r��C�K>����̞�[��5�崉6�w��}
�z�R�7����w���k'݋:컧�����J���-���E���J���@�+�(��x� !Қ�k��A��h���x�mb�׊�k����7Ζ�VOL�; �y�z��>���h\���&���Kb�����K�6���������?�ːO���Q�1&K���T��D�p/2�qu�n}d=�{��~�6���+�PP���g(�dF�)�#�>�> \ؖ�N��d��4�H�G��m!s�7A��H�����
v��K��38)�����R����}�!@͜`���au�xo�+��4�����P�0����@���?2�}�N��3iG;�ە!P�}��>��XKM
�$Vp��>�J�+��n�G�V3��1BR�O����`E�|�Qtd�8M��h�|X�j\�JZ]!�G���u��Y��x秺B'Ƙ�n\I��U�0l	t� ?��E�!�k�Ͼy�cd�\���wk����7��@����!�cB(��bb`x�Փ��FM!kܶ�2Ȝ����s~|�6�ο���sX�0h���^*k6e�����cM;Ґ�
VUȚ���ܥ�n�� ���b����,��*�f�hC�!����|$g1��,�e:.9]ez�i.��^-���{�jo��$����H.qR�o?�(M�2y��z�R�x��O��Qc�~����S��LNBd$��1~��7�;��d)�p�������{ E�A����(�R�b����R<��'/5��~������n/l�+�l��6�F�!��-"`/R]��b=�9�>g�Ç夷�q�����߫���i��Fa{�S�Kyyg�� �հ��Z�1�e�3�v�׵��(7D�z���yS��LM�_ǔ$��b��Kb��SW�.&�l���8���<�M������"�;��Na������ҋ-��h�Έ�|Ԏ���ۗZ)�	���Y��F��mdPʽ0T����.�m���܉?���)�f�nH��X����r�'�3�������/��__�?�ɢ$��T�$\1����<{Rq�4�:�$ń؜ �l�DL�aA��g�Z�&%����H����K�B���(�x$rVz�8>*ק��r�;]�L#�'���� �-bN�ت��s�(���DXyWH
%�Q�	ܕK�W:5�r��Dr��n��
����[^�����FX/C3a�3�hb0k�F���Y��W�s�0f?fa]�C���D���]�>��*rukzm1C�Q�W*K2�\��%"'\�����F�A�ڄHu1��Ԍ��O���ۍ��4���$��0fW������FrӶa�eB�"GC�i�Z�R8tC�_��}Ab<���ug��W!���}SV���w�P�"1��BB��Z��l�T�e
�D����p�h��C�>��Z�y�M���R+�1�(�tp�UE�
�@U�-�P�w�Z�} ��r�ϸn�r�q��n����9}��]������=l�ۧ���ӯ$��r�x�+�#�#d�E���ڻ�����vLs<K��Iؤ�v�ӡ���a��t��i��������W���������hm��#L|F�7�F��+5n4O��$���y�(p��,,�x�J���m\��5���	��# �J�dP���5{����|�� _�с#͏�����]
��y���{T!��R,p�a��w=�w�%���}#�L�S�T�V8��hzG��fFo=�G����*��^�S0����p���K.��	���(�"F�'���S��y�M�M�0_�I�P,h��x�����m���*��1��/�y�Y��XՔ���+�BR�*t�~��wLL�S3�����<�^Lpע���-��r]TZ�.hw��c��>�Z{�I�FY���/�!Nw��I�4G;��Z�J"���#|vO4�\�\��On1h�xE��9-�ŵ����v�"B��3'k�@1)�3E��ʞ�w֙����z��=�m6�ϒ����ӓ�=�l�UPՊ�O.�Zۛ����ݑ!��;�l�I*�v���0Ot�4�� �"G�bH�:2�3jE)�&��gQ���aM�ҝHء�RT�)$,'����m�V���
�hC�tѺ����g�%�2F�5�� ˔���Z}E�l.�5�>z� V���N�j���~2����~�Bo�� �ߍH�6����#Y�UOs�~)}T���`�6�$�;��߰��O�=��z�����%�d'�?u�i8�Ӓj�l�74Zq�5�'����ó��
���|�)#Y��p�F�w�H�����<C�_,÷����Ϝ��"_)����5��ǯ&��DZCUA�d6��öҧ&.g�.��b_.�.��6�7?(o*G��a��U�X/R�Tl�:��n:�J0����	������|�JT+�"�y��E�K�奸]nE�b�L~���}�8���:�C`0�mnaB�^�$���̜�ӣ3���k��̿; z���"��x����ήq�|�K�Ҍ��mc㉂���xTd�p4��t����E�S�(���&�	ϘMrҿ�d��q7������2	fY=)�2�k|f������P�6�D��	�(��Ɇ_H��b���j��yεz^�`�ĵ�΀�ߟw�B:9�ռS��=�����ug�2C���K����|��#熾�Q��GЙ}\AH�D�ɘ���)��־Kv�>���<-�0�܅=�@� 5�w|��\�yH��Z1��x���#;{@�Zp�o�li<��phT^��˞r�N3"��t�6�0� d�|C�'���r��f�3�K�n��%��Z��0�����`��c^�YK�����I�P������h1�90U��[�c:@n�oj���*dx0��!X��j�%�\t$��t�����q|>@�� �prGw���b�Pذ`|8�es�J��2�.R���\U�-#*�2$��~O��Z��F*�*��5�:�Jm�yA�ad��S��U��������d��E}v���K�K�%U�?��������l�G�����n�5>)��Ԍ'z%�J�pu^D�s�r��G���]�C�U��-%�R��H��Z�R��\~Bw?ێ>&�j�5}�t�k���+�̓x����#�IV�'��]	$7��"j�.=��䗒NXЉ�b LjѤ�Ɯ�)O��gz
M��W�A�,'�*�]���e�sw��("��I
TP���G;����)�Lg7�G��`xpM�0�?鶻��\dP��k-R�3*�ўgo��Y\3V4_)HB�b�O����7���B�[4/Y���M$Z�K���jf^J�8ވG�L��F<@L����rM�{����+���0�ykv�`E�rЀ�[��
w~��h��P$�ݼߕ�B��d'8(u�r��t�&�/��y�I�����|RA#�I��v^e㢪���}���_G���n��^)�0U�ë.�r,�u��q��[�ɒ�~�q��Qt�y𙞛d�q�������o���A��GkI����{P|D�:b:y��-����xS���6�A�@ꁔ�O��"+hm�����+N	���'�ԃ�_K�p(�����"�,���ֵ�e���e^�;�>n_W�����'�TN2�O�lt@�4��*����������mf��rT���_��J�u�5�XH*���� Pq��|��۽𡰽l4�@�����
�L� 7�y�  ��}B�O.^�eы֏v���)�+!��k|D��l�4��`*�ɥG���Ɂ��cQ娆(.B���p#"��z���ݵ(M�y���FL\��H��-�� ʴA�<:Bvϙ���{:?��U������?{!q��=�@שiWtNK ��gk"L�.����0Bj��?ez�ſi0lS��C��Y��*��srW�&��Λ�VvBe=����JG�txNЩ�`7l��j�$���U6�#�������˓Y���3 {��j_�E{�z�x��Fګ�6�Z�H�_�o�qg,�B<L�)F+��opA�*19�+z�����x7`cSmn�#"a2�3�j�~��v�
�(��$<k U�ߌ�4g��$��)�[&��V_q5J�O�|��{1 ��|�Ȇ2�������> ��O��Ls��f1D��\]
��ip0���v�_e|�L�R��-=+|i��|k9L����i�֯\�6g�g�<_�fKMC#���yR���m� ��)&_��G�I��S��:�fױ"ۙ�n��V�JI
�B͒�
Z'�=�'���=�Sd�`�����>>)�$ڲ}#g�_���q�%�٤���y;��?����a�鎹 �E}�*��L������p�ca�E�j4��5HS�*���;��߃�@��m�ꅾR�=y�񡡔o��3�����m�}Յ��� ���j��Gڃ�يג�YJ�n5Ia[���S|��B�#�����B�(��{R��6|8���+J����v[���^�v�IF��0x��Q�p�hc�s|�՗bZ������Q��
�2h��u��U6�k�PL��Z��1cŹb}5Y%R�)0����08k���s<�����B��T�����'�1�e�R��1�]�c��2ڤZ�n ��p1|V�@��@%8T�N�B:e�����kȧ����:��e�~�h��[L���4��\��b�PG`#W��!õW�ll�*�*�6 �!� �!B�W��գSS�徺֢m~�m���Q�e�3���*�[�*��E�Wp;ҍfU=l�<���nX��:"Q8{�(>X���j��b�������ɻ��hQ����b{��)���&4s��R9�ԗ��u�h?�?o����&}���]8���/�!VA�������9�瓣6�)s�z�Np���(�[�ê�HЈ�&���l100�uN;�%�+b̐'̞ƀɍSb�>�!}%�9��+�j��ZB�=b�1��ub�#�R0��5ur��Jv�Q����F�9Fx�jq�:��Bz_k��p�����F������K�m�^<M����w��)E~��.��{ؿ{�u��MJUT��wfێ=��3p�������G�ϑ6-'p�����3gF�,u����'�p_ 1�����SB*�۞�A�a����$#��J����"c (�s�ʄSv1�8s9�C�$���M}��
���ъ�z�u�/�ĩ�w��P@<�'y�3ں��
[��&�ӔA"ڌ������_�ױjy6V�) I+��!��P��rIU���RMbR���;
LMrv�]x��6��\��"yڂ$�逖!jz�}:���exZ8���F_@��*+Z�U�t1�сrk � �ֲ�r�/|m�K>6�>R[�37�vA�e�KAp���v��_��[t��p���M�c�΂?�����[L��(��0Z��W�j��|���Z������󟍘�Ɍ*G�Q��'�~��!`�Y7����{R��\�|%��d/"��36���`4�i��h�D�u%���
��L0���2Cх�v(^�2�Y<J��ʨ^�\b��%H�h-�����-R2���N�=��|�� �b��X0��ɌS0�Aق�)j�������i��p�RW�+�Z��{p!���<u�l��:'T�TfY�*]&]&�7ः,A�Xx��rQIX��?H�4������Ys��Il�yXc�7U�����3&S�+j�����PG���a��{�e�,vj��n�����b���d��if@?�"���>Pw���2k����r�r�;
��F~�����W����3��� R�k�;�Q�G�
[�A�{��yぉ&���T��~䵇��i�_�r��%d�s9t��B;����W�"_�j�*�K��*Bc}|���b��u�o~Q��~��l�;� p��,���7��sDL�dz����k��x�Ƥ4��6)����jX
����oI�+/�=��ӌQ� �>Ax��n3rl0T��r�	H��OB$�џ/�z�y��r`	��r0.-疙�߿h�߯���O}
�U˙GG8��y�O�?�,�0�4_蔘�'e m�7�W�?X4�o����p�xTd�{n�l�4���Qɴ�����n�t6=�-��\��������ԎCȬ�VO�tr���c�3�})���3"(��:>���u�~��%����!�^>8��z����r�3�d��½����^�>8	�hP�"�I%�Jѡ��c�	N
�F�O��oS��'�q6s�v���Z�-�c ��,;��S�WH>+jBX��q�ד/��A��²���ќy���Kd2H��T�Ψٰ_���VE�P����O�̣ծ̏���i
�ֿW��X���5LC��ږ�����E��o�5�Y�Bx���.1�{�:�̉�e�qc�b-k�n"�M�r�)Gm�w65c.�@m�1���hKW]���<��R�HfD����KաHS�7���~��<���q[����Ry,�|8�LW���Jf��J9��Z�u�Z@�\M��"#Z}��;)aT6�KJH\
')pe�lZ
a�f�y��(��?��k�3B�O����I"OWu��L��$��H}�L�ߚ"��(�S���� �GAm�����e��4�m����,�'��M��+D�d*�(���8!Pq�V�'\�[�9��
�kF0᧚dA]��p^h0��vϱk�隺w/�d$Q_/���
l�J" �@��Ы;���H���e�C@9	q2&اK�����}���� ��X�,��Ys���0)k+�Gլ ���L�xpa�5a ��6�M~1��H�V(������
^�XK�INE�+��V�6E�qn%���F��W�y���k�"]�c��_t��c3�
�o�\�J3ZI����	�1��eаeRȐ{U��ٔ\5h����jP)��uӨ:�p0�pNa�UǮ�,8Z�*��M��]S�:������v=�Sց��$r��Tc�a2+MjwwK���I6�~�a=Z�_!&����VZ���	-X���Kf�A�H%�Ql��ȃ�e�S�.H��}Q#��2ٮ�_eK�݅��E�anWxM�j��*�^Q`_TjUy9i�r�/9��6��L�^�x��cH�x��sj������޸u�u�Pj!ѵvLN_�RgR��{m�{���Ղʢ��s�3R^��USF�Kn�SLK�`�`���uz�_;,�BY��;����b�e����`�-9�زr�8��8�moQ�/p��l_G�X�na�����
�ȥ�v9�����E�b�>���L������,��P�@M.��#_
�w{����P
���6�:�X> ߇Mk#��}��|��ئ2 ~�6v� �y8f�otx�g'uV�=uH�,��ރ<�n���F��<g��Xوi�[C�A�<�481_�)��#��v��TS+���A���2z�$.���?L1���,I����j��Z俍�g���&ow�>w3~v)-f�g.{��z�ݨ��ÀF�x��z1/r�)G���*�����&§	�[2�`��t��>�5��܃�j\b�`�fI�4����e�[����"�G���N��3{ZUk��gM|�'�t#O̲e�k���2(	����2�D�<��v�4�Zb����h��մa�rqC?0Bx��e��M�n��l�5��vr	���m��u�z��i���O�@�L�E��C�/$���K��-��=g�,6�@!s��
�um��9��B^O�q������n�^��;��2���<8�����S:�f�vc3M6���m�.;K��R^W�p����q8�l�A��� �C
��nJ�&�E�N����"�J^�K�`�D�� ���GE���I��\5��&��|�IsXZ�a(�v��N��<,ܳE*|k,���/�ߨL�`g���g'��e�^�r�LC��R#�U�:OR����l������qrH�����J%l��\]t�)�6�Il{��n='sy��f
����ۑȳS����C�(Z�+N��"I�-cǀ�CQ�YV�}�ȡ��ɔ��m�g���4��8���O�*ђ&���z|��AK�[�:G������i�g!S�@E����:�`�����ܬ1fLX�F#�Ɨ�Y�3���*�B��9>r�&@x9�e�xߏv�7|����,fp�CJ=��)J����XC
�K�x/JWRx.�W�l�o-�gA�fw�=(вكl�2��>q\A��K�ce,}Xq���#ߨ��(�TM�\� �7����T_��m��]Liʭ85���/|O*���Ŧ�Qo�����VV�(U��k�u�u=@N��������_�~��+�v�e���W���t���>��G��{����8�)u�cD�������=���CLK�>)�ո%S�^���`�����Sa�4��^�56E,g��	&�DC�@��s�I)16wP�~�t��>~��/̑C��vZ��n�橴Gͦf�t&���vŔ@bp<2�����(��o&Oe .ɤz��f[�A���5d���>�ʂՂ�F ��~_7پ�}3W��}� ���ZPd{>���T�b}l�J�!��Ώ�k;՗�����~�J�z����O��~�0���<Gb��/DH��mp��o���t�c�F�vSc��b��(/xY+M��ny��$8�%0� 5������4�JR�TTs���1����x��<&ZhM�D?B����e�>:_4�d���iNE�g�QFN����Z�2���qy7��(���j��G�����,�L5!�%FP��p.\
[�����r�Ѥ_"W���܀6z�K����^R�Mm�]��h橔 F�x�B,�Ј��mt5��YXd�D8>K�0׋�5�Y�i�B��ų�= ��o7U\�1y��!�Eu���~������*-biyt�`����:�}X��e7����:τ�j��$b�j?�j��`�j��.��j}U��Y�Bߍ�]n	w�c	e}HA��_Sِ�8$�82�C�5І(�_DU�"� ��ȭ-�eqZY��MŢ�֪D6���J|�^��+Q��;���p�UZ�&+rEe��> ��Jm��1$f����nb��.�&���vɩ���z�c-ݾ��k��o��ؗ�ĵ��5��(�����䗲O���(hZo���6߃����M�&v:#{��.XR0<�z�{�Μ�\ШK�{e���'F��]��4aQ�0*p9tp�$l�ez�l/�lI1���!%�31_J2\h���J�|aXkKG%�#��M��סG`�\���@w�����H�M(���\bCx�e�.�Ě�Oh�k���4�I�`rq�a�i.��J�]l�+z�k,]gWORm�<�2 ��TVz��ހ�ҥ��`�Z%Ҧȼtv� *����S����
T=��H���OG;�_ܜ �K!{��q�㡇�smҝ�,+0n���L�:��x�"���<�5 �/#��٭rJ�Q��k^��.���=�l���ĻTċ!��.P�t�v=��������6���D�r�V�$��b�W�=C��q�(��s�������6p��-����Q�+NM^)�~6.l,�-��³�ÞA�p��4q㟉4g&� W�jA^mP}~a�g��BLkE֣�6@xV�u��c�4>���(�|�"x��V�J�􁳓0ē�/��
�QO�<�_�M��|��ƻ���C��gR'b%�or�Ka��՞jRpO�ճ���=ª�%v
�%���i�����ſlj+�z��2/��ZK���������S��bZ�{A���L���̪�s�T�C�s'
"��)Kk3΃x@U��xww��}f�
�DvO� -�˯�mȣ�H�σ:��ۭB�W�D���߬򇃾�7���7h�M:_k�������^"�2ã��(���	�{�3T>��t/Y<�)&�5L���~�4̲%�Plh����]��e+�btM�8cI1h����{�
B�t��Jd�}t4eC.��@Q��R�*Q��FC�b��>n���Y8L
��`Vg>�b���`���?)��Cn�����D�rQ��T����`�B��������Z#=>\$���9�gn��북jǔH����M���'X��o�*l��]4��h��Bb$�*%�{#L�dӮ��䪱1y�|��#A�ٵ8^���Ӄ�l�k�k��m	����(���^䄝v/��&��) ����l����s-gS�bbҶ�-�p�R%p�WJŚ6� �j�2�sw6��� �$~|��PP�Pq���sU*���@Uݡ�8�W,�&�5+���֠)����֮����я�X�E1:g�Jߟ���J�A�)n!|4u����;X+jn(�;C	�d7�;��|��9�o�A��! �3� ����j�)E2��l���L9+��9R=����H]2:��ӈCi���y|O�8�{R�M����}R����$#�F��0���5SV�Ɣ�1E�
��I�b�gp
*ԃ�V|��*z�z��5�i�D�A�zT&vO���͍+ɖ����d��-yh�|P����𕣓�Z�wv��B�J�4o�N|C���b5��0	?W��#1�`=)���'�u��������'U`	�FO�X���Yl����K`�+�ػ࿼�rM{�HYFw��҂�'I�]�z�Rݡ��~H����x�os�c��Κ�є�ȓ}��|^OC�V��UL�P�����+°�_�^��Io�$C��zBҟPo�6|P����9���1�t��;}a\�gv$ʍݱܕ
s�x���tL�Rpl$�Q���[��;`���ʗg^1��#���Z�h�όj
�~���t�D�L^)f��E��U������JZk�X�V
G]g�A��GT��p48�~������ɽfrAN�a���ԕ���1YҘ�|xG���/m/������1�JƔ􀺧~�֝��dr"�����%t���w]/oB(�F1�g��N��*�J�0�k��$ �S�uPM��Q�a�v�����g����
�0l4<�Hb%

_j�d�u��xx6�R��L&X�=��L�;���O~�ګ�A�}^<����Gv�|&2��\����l��kS|�k�u���R>}��;]����M��o�fp6�i������������3��Zjsә���'^��6K�GB��S��� ;��Z���dG�B2���A���i>#�oJ�ؙ%�Eϛ���/*A��YvQ�Kv����^�qŮ�X֔�bW<�6* �L6�^�y4cv�0��)���f�T���r�e�~�e�}�3{+@r?�g��bb5>0��NWPVQ���n�B�(I�3���<+�~e����#�ǀ�z��V�P�VP�q`�n��o�������,����jf���\i�V+�=���$@��s��M*�e�'3�5�#�<�0��6i�7��m,�h�?1y��C�T��:�
r�� 2�B�g�d�W)��%C���3br��_ej��C�4U �Ɠ#���V'��mT=�;}/�i:B���joB�v?�]pJ�x˩U�5T���GqM-9�� ��Ѿ���Y|���&��RZ��]8�nv��B�+E�<u����Rp�R6���,�2�W�T����=?�&���MVK�qǵ��IQc�,S����+Xz5!~��HF=@�WO�{�Q������)Y��Ee�n�_N�6�p�oo3�6Pr꿕�3:��~��a�?�z}���K{�(�Be��D��k[g�)졩/
�O�!��p\ˣ�S���I�l��]k=qM���b�I�_ov�F��#����qrm����0���Mo���Vq��'b�ȿ�J(���u�$��K��v$��	 ŏ�Ӿ$�O`�h4�F��I���G�p��J'49q�ue<�9B�g�D��JO�#9"�}���Izsb���$^���Se��m(�	���q�E?�$�9(\B򎺪F�Ӽ/�M����%�*tuݑ1��`��N�*��n�!q��rR�>g	���8 4-�Ӛ��u�� ]�Ѱ"�ΧR��	�l��<L�L�"���\�?&����9�
O�N�o#V�4T�mV�mHб���F6C@�W0/��_v3��{�~#Z&�Bb�2�S;e��u�����z�3���b9�1<U�6AJ��Ҋ����j�W\�C��p�f(�{٨���Aν������G(? ��5�4f��"����*�}�j;	?��7]2c
Ј��n� ��{/�C�Ί\.)�~��� ���"�V�� #�W+h �cB�5`��v���<��ڀ5�C0�|��*����������a��	A8��0�T8>Nj��S�s�
������,�fA��s�Ѯ9O�+�'i�"���`�������d�8�E�ߙ �ۜ���G`g���Ü@T�$֪�>���ID7��JD��F��[�髋B�,|T���g��	Y9�c��,&�0�x8R5Z�><�?T��^:K��I~�?B�����k`���9�� '�\�U��`����D���::�]��k����G=�j�0��#�]m���K W3�W�-��U��f&Ϣ�L��P�/!�S;JD�����]EBnF��Q#�#��jý�JxO�>�a�,0
��yJg�O\w��(��2�lˆ1�{���+;HO�vb=_���N��P�Α�|u!��Auˎy:H ��+���<T�� Gw�姥C�˄^�C)��f���2�
 dX�� ��s�N�媝�gF���)��q]k-vB/�-�s6ۢ1()*	��0�TT�EMҲ��F�g�kw�$7����w�7�0|Y폾�WwqBY���"8ZKo�OR)d��lvv�����r�ڜ��َ*���,D��&+�L�e|�!��Y�zI(ej�):��EG^OJ�9cn���8�I�7��kj��w�.��{���8sg$9T9:^&H�D�5T*u��Ή/�����i !CA%�-^S��I)J#,Q�0�?�I��;.&��4����9���&.0,:�
m���̸`_�
�n _�º���c5xatC��j؊��#kWۊ��������/�d�:���2�cb]sC-y���e�*8�$�Eɿ��`"M�qY�8=����_�[!y���ô9|to���A&>���sµ9(����G�r��[f,�
B�x�F]�^�~��J��;E3�{e���[�#�R�i�`d��nD:G�O��P��Cu��v]��)��]*��F���Wx�@�4K�?�<�!�h�J.|VFɢs�(�i����ϦW��Js���H��`����x��:Ǻ|�^ƛkyA�/ !q���g�-q,Bg��ҹΙ.�M�Kc�*G,A���LFD��OL�ܢ�����mKC�s&�p���Y�	�	i�:'��sZ�ۺ���Ō6��Ԋp��J�ʼ��j��
H�/Ꙕ�h82_f�R��y�1�'����D�(F�N�d�ӍF�j[��C�U���C@y�����	�\�}��,�%���N������`�7K*��/��B�%z�W*-\6�ֈ���J�`�W�&�.s��e�WzF�uW�rEda�ܜ	J��pa�k`R��V��8l?�
��d#�d�y���$|��W�p?<+��(���K`0��X{�	M�߀t���^�%}�X��/�1r{DŁ��KK]����GZ�J":E�fC7�Ӽ#��P���n�
a.#�B�����rO4cȪw���y�/&'�#�Ӣ�	�7 ?ڡ��{\�'�&<��R��&�e�x)h8�	�B.r��w��Ґ~�F�x��(
UB$�n0�as���S�x��@X���C����?��ǩ��j�6�*���=�L'T�V�]!��VKD* &�3rT����AT��LFD8��oS4��c�e|3q�!��e�_yZ$L6�ྎK�}�t>�g�Ǉ��N��i�`���P������J�^�g��� ڛK��~��3,�$�ڹ;T�b�r6#N՛�z���~>�l�����b����>�vڋ�*'9���^�P�7�����$���q������fxF2Gn�����Iĭ)]���~*BH��I]5�p����nP��Qn5sJ�6�-��*#6z���U��Ͽ�VHi\�rqV�+�A���b+�����Xc17KÖ �σW�]���K�ګАj�sn`�Lp]�>�����Ú��]���b8���H{*ī�8S�>�|%�B7)�����������S<zg����ܠ��y@�Eb����錄�"5��,�o!�����a�\�/Q�Ft�
G���wDN��x�udy:>b�g	|AD�A:ms��l��A�$S���¸��刭��)�sM�ɒ;�O��,ԗ�1?#N�)��a��H[l�a����?S b�B�Oe^�����8�3:��b�����������#��k&�˯t,?G������������V)7��]^�|0s
� C�����a� z��)��=(���区�?i؏�O"��o��Kƌm���h/�=����6�����+��D�[Vc�.�b�ҕ�*�F���-p����2����*��ۧ`~�.�1��<��nzE7�mҾ���E
�FPF��5��]lo�ꪣ;ՈM9�U��	^.��n��GBU�`'<[���*���WL�h 8R��y��F0����|��룁D�
%��)�_�	�ꕚfM�h0�n�5k`���|����fD�u5�w����H7�N���<lµ �1_��V�xY����2(�����b�!�� ��%2p3K�4��3�q���'l� ,��upnu#I����z�w���`Ƙ�3��&=b�g�;y2��삹w��P���j������]Y�\�RV�pXJ`2<Һ���:
m�L�w4pO�Yoyuk�<@øvp�L�5E5:P��o_�R�����1�ϲ	鞜N�S�W�4C�1H^j��*�ҿ7�# ��"���zY��u-��6��;b=���"�P��@���9�6�;_X��T�?��a����z��#5Oj�+�W�_^Ɛ3#sؠ�����&j �UW�3��ɘ�%1��J�����֨L>N��}昅d<p{�2���Q���#�$�ΰ�QC�(���5ֹ�c��y��r��0����� �MIВ�rǚp2���S� ^��8�� <����CqC��ʂLSc�.�x�)x�}�����R�,�1�	���zU����	�bu�bL�k�ewPs�g(x���:[:q�L@��)�BH���{���;cCa��P�^o����T��,�gu<�*�u/�ƺՏ��4摧��z���>7�g������E�͹6�����zw���K3�A���C݊�t�x���:��O'�ҳ]+ICS�������d~�
Z��;D�K�\�HU������;�j�n*�<6Y�Z�)F}h�R6��D2�-zx�Wo1n�>J�_��y�w8�����l��.�5��{b'�Ս$��U�3C%KI;�l��K��3^��m*]Ʒi2���X�&���d#�e��o������NB�d+-*��('y#��M�Ҽ*��N%�\���$I8�P$����3�O��Y�>�|�@��(t p�t�;�J�ٜyzG�M��r�>��Z����&%���b ~tK�h|7wh)��X7�����W��<��@���
l�qf#I,@�V�S�0�+��cJ"��ץN#0,(�Wk����{TQ��5y���Έ���j!q`u�<� V���%��Z��V|�P���c�"��.Yc�>Gb=�	�+��ߣƚٲ Joj��!�Q����h�o�=:�K��T1��VH6�����oY�9����!#��jdjN����i���}�	.3M�F���PLQ���UĹCu&�=�=#6�~c�\�����կ��b1;r<�6��JzؓQ�gdK��*菔I� �_��Q�7sj��~�^��tu?��F	�=��E�����첥_N�d���A��[�l�0�/D��ZDA�(��c�)��d�+E��o� �K�U`��?�8~4)�J�)����h�THv�z[���B�۱�C~�ТN��~�v�1�$�C%�����#:��N�ONM��ϔ}zީ��z��B]���$��cSa�5l���0��
IwԐ�����*�i�<y^R��v��1��6�>�U������)S^9��y�{��
���CLUU�1}kb�6������=@U�~�/��a�"�Mr�f��z�[�d��:�E�vq��T�NE=X�DP&��a>Yzn�|G�Y��ZB畭�o�+=t�Q��.��l�`��{���jv{~���&�#����;ɗҁ+��B�>�	��|Z7���lT��~tDB.	*�+�'�A���ul}��P�w��i=���e+�ܝu�G%���F�:�vN�Dӥ`l*Mr����q��e��j!�G�ٸ�Oc�hϘ�Z��F�y�ǇG�%i:@��j�M�ԗ�;Q�zR(�qq_��v��K�G��C�Q�<E Ǜ�,.����,U+�+$X(C�,�_)��+z�/V�gbp.�=H�\�0������j�9��܃MM��X����~w��N���`��_1	�0�3w��V��9M����mnP*�V:	�r���w�.v�����a�Ee�	�Ns�|� .z�Q]<�{����qr��L5�T򲅂�Ў�h|͕k�ة�Λc-�O�g%�{�聛VF�)���u�-&M��@R��?ji�<�mJ�qmՄ�FL�~���*�Aub���A�D,����>��T���"������Q��8W�L��IC��k���I~��EUb��� ��2$Ͼ�~��3���kP����`1
<���9H���L#sU�������q ���Lj���o�8c��~�[)��H�\|pV�m>��+�o�7���{��&P{�/����eU�����u(�?=��حB:�%���f�-^�g�������@�:B�(�L�{����Dى�`��;FC�:�9Ƙ��M_4_��3�&�ύ<\@i�q���O����� �J�K�7j�W���S�7n��}����ŶCwo��d�'6�HO�;�ȣ�Q�w5E��i�J�#1��R�ݠSX ��c�����j�>\޳o�����kS����g!ZW�l�o�h��Q�1����K��X�t��bF��u�dV�DKjazb�ƕ|g1�$5p>y=�s% ���1Dt��T�B��6ޗ\
`���e����`rÅBR�O֣8�+i�j������E�?�Ў�fv/��?��[��07���W�_��@f�%b���Wc�t1{nƩI}��	WE�&��J��,x�r����Y8ڍ;W)��� �%��ھ�-��`w/lǝh��e=��\zB"^�[:7`�%���l>J���� KEw�@H��׆��>�3�F��a?�ċB�lt:�N�����q����Z��*P�������7Wl���S]�"��*
�&qo��:'.�Q��ftU�i�x5��V�w
����B 9�%���~��.���a�X�H�|CӍk�������.��|�=��d����g.��,�����M�s��XF+�R�v��{�qwz��s��I�
z��q+�l���������'*���}KR�)�F�D��V�8w��{1xV؝��ev�|5��P<�ͣ1+*<���F|z�H���M�>qǞh��r
�\����� +���&���#����J[�?:I��So!D��Q�0n��;*�q�{K+���;��N)�T�T<D�D�Bp ᴓ�ҙ���Di#���T��GR��f����x��8�����E{����u k3A�>�7�Z�����E�FL�;6X��Հ���s¦�\{�#,���V�������j��:�y[5807:N#��E�"�,�#-d�'�/��BH�/lU-%�������T d1t��]$�9^Խ���r��:<B��e���G�����I�C�[�I��O�z�E���%�&@CR1�E����s��kӄ� ��/Ų�?�Zר��o�	�f��G��|����Ez�ې��'z��m7q�h�IR&� DQP����"muTAk#�2pD�[QE��T�	}�î�2/B��ʬ"�z����_�W~/�.r�g���F���  
���F�(	�6����'#��xMZ�c	dI�uTV���c�7p�_1�R��GT����ֽD-ΊET;�'aUFW���,�S���5�'�G��9̔��1-.Ø�MS��(�ʲ���^�`N����Ǐ^�{��O�7.���#�$6!�V�#��/l�~. ���=)��� f2°*�&�K8[g4*m����]󛫸iv6�~ήүa]�1��8�	ޜ���L�51QI�L�31_Yl�
$rM�K��c��4Hıs�{�J����U����^@�����Hjy�6�����
�N��,=�nq��~C����z����_�#��)�_&OvR�������������_�^��G}vCn5�8z�5e�,@�E�g�Mw��t4p��KLP��q��Y����
�7�p:�
a�Ә/���F��Aօ��ͽ-����RZ7K�l�ћ�>��)�oQk�G���}��nv#�4ƴɓ5��`1�Go) �D�GޘT�due(��J�<�
YdI��&�l�1,�<���'����m���%i�GsK������y���ԚT)O����sĪ}l� y[�5��Y�O�L�R�HOU��k0q����}���=Ef:��q��l~׮s^�r��/�k3�5|{q��/�����.�����)Yq�G����.ymZUY�QU�ms�(s������U�6�sb���!�_�z�z�[��D� ~�������f2~�1�(��
��+�/f~6�"��X]�h�Q����Y�����I�ؾI���K�˲dp{f�D�w�*��:�{~�`� o��i"�c��`���s����	�4:P�=:0�n�M41���S������Z�0�
@�=%&��\>�~<s��-yh����<�w?X�^�=���U��fa�AS�m�aE���4?��{��E�.t�cӥ��otB��	"�Բc po6oN'N��d KQV�K��d���}Y(t��;��R����gy��7�#Qsб���.o�˲�S��@!_Z�Kx�7����>�% ._q8%��Un�:dOc���s���cOx��߼�:�����o�,��f+�c#�%ESjTzn���Plªe�.�/}<Z�u8m.��f�!j"�3�Ep�8��}���Z"�Hq`�0_M\:�:���X��ChR�R�1=]X����93�&Оd�2�"jc�̅"%�$_nߚ�vh\Д<�N��s�wPD�Y��eu�M�L\3�%ꇂ��=�[eߞt�JM6Yy��ulo� ��B��l�
_	�������Qn?<LX��/����B��\����$��i��g����/-�M�"c�E�vH_f�q܉$��$1Nr�~�;�n��d*ği��R�U福�M�U�\z��ypB�i�Ŭ����A40�ȲL\M���׃��7�ʌn�Kc�|,�P�l�i��x;qŕ��V����Y�9\yt�1 �e擅����I<��u^Gy�l!S$�P��*��J�AdGk�a����A�$=h�]�}��KynhWrJ{�y�b|��PG�xM�K�h~@~�Z��3��Sӷ�L��e)F&�,�۩�	ϊ(uH�R�,���=@��Y��|�.Ak�Ӌ~�ُKL��M�h�9��I�cZ�Gۮ�覕���e-��o�F@*-N]��	�3b,��Kʡ�Y�6�q��ޗ],B}�k(:�����"8�DF����&��no�A�[�+MW�|�6e�,�H�m����E�/\�+�{�:�
[�Q��cJ��_�;������7��h�E3�<��C9�⯁�K��٢�q�j�m��R_���G�2��7�ݚ������ܤ��?����S3�Տ����#�k�7:v9@�G���1���B|0Ҿ�i\�� �'}RN��c�9����i�V��o1K�&O>�Y���C�����r2��X���fj��L޶�s��]T���ʹ��L�����n��l��B(}�s�E%:����:��<]�~æ���>_x穈6��(?���	�"��H=��n��A1��ޔ��E��a'�)�����Ϳ�W�wG��[� GW�"�;X	����l���U�r��8�J	�w"��+hzTI��lQ�j��?�[[�Ȑ�%����w٭���#�u2/I�Ӕ�(&��Ҋy$x��+NG��F* ��:�ֻ���Δ�6'��3W׽O�*/,����6$e�F��a����Þ�6֋n��l��v�=.�HJ���
7u����CE�M(�'I6"�m�Ax�'|��QJ�]H��7:f5����J�϶Xs�?�6 ���7���w}�7���e���:��|���=�#�+_�o�Y*v���l`X5$l7��F�i��$ă`\u�-"@s��]wX���coX$�~uX��������y��#��b��oˌ��
�C/��v�r�
Fqx8��b�w�͞���N��� �����34�cU�K6gʄ�w
�,̦�����gޒ'�8���}�vf����K�|����q��§���:��?w-����]X<�07�M�q��0wC��tJb��L������=?X�6/6���f̫��յ5s߱Li �ƺ���|��`�	t�j+��-8#J�����d�.��;_����޶4�����\Ԡ��y��J&�׬��K��t�ˣ[-<t,Jz�mG��ჳ^b5p9A���\��!<~�o�� �,��含G`O"��� �.��A��s��L�Ԍ�=B�����>�{��F��)�@0F�NU��}�D����)x��L-�21����,?�w��ų.��ڰ�(�0I~���о_{,��5������� �V�'~"j{~��S�@��4�R5_7Żt5�DXW�cƶ8����V�ō���)��#�lϕP��-��xB��uu�z�%Yۉ㥋V���Ѓsk�ʹ���Z������<��v+m��t�4��"���(c���F��94�|@6��W�+0u-�Q/���&�$�#Y��O��q��y���:-�0����047e�*��+C�vG[���:F��FVBwu�iL�e}؝ぉ%R$��F6� x�(��P���D��B>�(dPP!-��;�����'S �z��c��������b���1�f�{�[yOgK1
9�2�_�i�ͣ:b��rSğؔZ�Pf��8�K,S�z�fxA�%��<��X�Aئ��J��̢��X���Ӭ3�Л86�p ���e�ɓ6�iǸ<M�X� @�Go��'���;J�T�e�XtfeJ-�z9�{�Z�k(�X����a�� ������}oޥ
��9/��^�K\|�Ţ1/`�a�>K�/�odu�B���*����:f�D�&{l5����v��L���a^� �)!��0%<�ejzp��ԍ��k�c����z�߉�2\���e"k�wF��B�e���_Lҷ��~��ɥ��eӿ��D:_��A �p`�೜	�>���[}�p�v&Oz.��\�/N�k�������1��L`�����Q.i��pR��� L0`>�~"���zf�V�H�E4c>4��\x5`��w��))��)�����ڕ���Z�[Q 1ڄ��NI�ěN�OIu����XH���@����1��%8�:x���G�%��$k2�y�V`'m� (��j���v\�n��mR���q�����:�����yFC����g��o��w�
��Q�Ŧ̐l����cwC�l�o^�����`�������P��a��c�� e�m�r�������đ*�2��0va�.2r�
eE���۴�;�x��Z�u�ݨ	��u��½��8?=��ۋ��Q�Ie�^��ٮ��ƛ����-4�"�i�6��}Q��$�Y�ł�����n��o��
��yu�<�;�r�q�͎�2�|��D#��V+s�Xx�?Վ��H�3�|hI�]/m r��Ȧ�m��Z=.Y�4�=�n�y�X;kJSʓ7Ɖ���hk�TERz��w��=���k�bAg�nG�B9��؎�_����x><d�!vW�k���2����E�*ʠǱ{+�������>�߬��K�QY���ԗدQL�!�U��"�j�_�DV����Ж�|��e�;���¥�d�G���`���t��H�{��:�Ӌ�����H�Z,g�]��	�Q�8uۚ�k{)z�y,�n?h	=a����5@��r�sc��ʜإ4�@�h�è�&L�9�og��7V��ǻǘ ��ڏ�LË�QP��ι�IbF(�|��4`�`v�˴��4:/���K�B/!�D;�l���CG��K"�f��2kOf<<��s��+/҉J����b.\��t��؏�W�v�$��.�#�@����O�_8�G���{|�Ko���<|v[6V�,xp���/����e�Xw�d���<cQ۳��zm�}~*�eK�B�]�0�|�I�"X�O%r����@�5/�R���<PC��K��~=�kAW��X�!�������3j�dV}��U�>A�)�%%\��Bu�������<P��������"|�ȧ8�tA�]��Q*����L��L
I�jቬ
�e��g��#ZҎ.�^�Z���=N��o���<2�ӈ�≳�f+RIWW �咁eG����4���, l���yJn�BɶGݐL�s<2^��D��?|z�.;'ՀJ�GN�7<�-Wm:vW��K��+�N5f�X������|OŇ�J�'�0�!�!�I�d�>��1�&^����O�
���P�������@�a@����;����^oaRգ��KB�L(c����뒪ߕ�be�V�gu��Q�XM��CD&d�����UdM� c��� �y5輦&B������U�θJt�R�"R�SZ���x��#='���X��R�qS[~]yݥ/�K���G홭zo�7��Ȋa�Y�=��z]Ν@�8�	F`�#���jp/�e�q!Cο5��A͵B�L�QXA&#ӯ���Ԇd�+��(RL���ss��耢��yf��W� υ�����J��P�lgg&�Q6�ѳ����a�d�7�[TN���{���Tl�����/�04�;ۍxhw#��C2�����yQ3XA�c�EST���6p;5Ej�0���0�W�T[?����g�$�U���Vt�C��[	.�˚@�?8���Ǵأ��x�����U�1B��[i�	j�ͬ�+��-�����U�Vdb�Yz��ռG����&ol��Ri<��{���)����:Z/B>�NzIѡ�c�J��9�ұ��T	��[��J�r�dB$6�l�	�]3 ��T?��y�t\E~��᦬���DQ.:֍d��<S[�����R/�uK!�l�a����5F�7}��?X�l#�_�߂�&AXh�O˻��Q]L0/|p�>�}�"+���Vի��mYuD���	'�GYl^��9L抐��lQ�Z�" g_V-�@�FD�ʐ?�qÆ�2~`^���D�a"����^kNDx�kAi�;��&t�n���K #�0��AO��E�oi(�5�Q��2ߧ���L��9!D�P�R�2%*O��z�$q��AL��U뻺\�`�ᗜ��ԗ,>�����&�lࠤ}�m��V� ���˄M0��!���������ᘰ���S�1�ݑlw��r/T����8���f� Z]��j
a�h��@E���K��b&=`[�F��� N��5�E�LLx��P��w5�*n7�q2��L�F��Nx�n&�B%_7s�LL^~�:��g�q�@���s�Q[(����\�C��6��9�0���.�����[�@{*� ����G�-�"�l.�h��%|P�H������^�E�ak��$J�0}Ӧ����Rʡ�P�ȌM�j"��>������̖�|�r.� 4˧���,>�t\�*yE�L3��:��Yt�~B���E"�bCT�&�-]�=I�7K��;W<aL���6�n�ƌ �;�1;�#�x�	�!��DS��l{r!����7m�J"ΔC��iӿy"����*t���[��Q��}oŊd�ѩ�L�<G�4�"�2#[X�E����? 2�o ow��3�OT����"�.Q�S$��wA[0�S���d�8O�r�z|e�ӛh]�
�|2�^Cx�Ӥ�)e���"y��)�I l�d��f�	��יW̴��UبM��Wn�`����t���ܿ��C���j�* ���O\�S@h�H=�T�$ ���gN��Az��4���uW��K	���t�~��] ���sy�4Ң���Y��$�~G��S�P������^�Te\�Vˡҍڵ��g�V�R̨1�s:�����H�M�S�c��Ū�Y��H/��*[��H�'�N���m�J��7���s'� Wi��2�;4w�	bs����<���A���1#�N�br$��\7�*w�Ρ<�
,{uT˔)�}ڝ���Jpk�櫼۔5k�!q�i������Z��$�k8����T�><�r�kH���@�M�+a�k����0�xp	P�6��4:�B����d�'��#�69Z���2�6��mv�G9�����KK�l��	^��)�%��'���`^B!���t� X�'�񙢽�ߦr���8g��.6c��?<N��,�x6��"8�-�p�[�<��Rf]�ӉԎ� ��Zx@]£8c�r@I����.9>"g���#��=�懏)ڧn��+��/�����f5�r�S����;Y��Z��m��NU��d��������������i'���l7m$�֦��p���+�Q�ƞ��`�#_�/�:��������v��
���Q'j�!=6��j�U��u}U�I1{r9���&���3�G��Ϊ�u�~=G��tw��\�~��Uw���"���[����`ȏ��2�/��ڐK���/\������qh����O/�7��.�р.i��iD$����Cn�'9�;`�N��W듦����<���$��,P��x���B��w����dY���+e��qUXg��}Vc��iܿ�?�ژ�a�Mg .Xh3��M`�th�����8�ǚY�_\��3��<�ϧ�d�0���Cs@�-����io+�����1�^���Dd� ��M"��9�3�Zt�|&ާC4�G����E?6i ��-�5���4��;����^�����.�JJ��¸��*�RzH���H}���z�t|��Q�_q���Փ��n�^u�Ǩj��SR�$Ǔ��bZ=7wU�vqZ��(�U��b�ڔ�:Y^��\_��z$VotZ�Y:��Ȫ�̲\&���cAp{Џ� 4a���9��NA�S�6p3(J�bl����v�ʵ!��_�9Hk& �Oqꇻ�=e_q	%�i�H���%�L���c��i��9NS�Ŋ�%�hj���W�,�� <|���)�w�8q�聨�'�l0(�X���Դ2��L<��ID5�&�k�3�����j��fM�H�2+w�%���uP��?.��~�q%h3���<�H��
�yB`�.o�gY"t���X�a�/u�v�/��N��N!ڃ�m�����@s/ŝAcY����2�%X@"֊�Fy�K���d�-v�E�& 3|�-�_�K��ZF8N+ߐf.�K#��=���v��mh��/�x[���@Dk٘�� w���'�����ȍD�0ߔ'����(KyM�z��e|3p�QJ4�~�~?�J���M��[�����m���C��ܭ�K-&�/��c��ɶ9���k��c�tHT�9 ԹCW�,���H�D�*�Oy�=	}��5�M!I�L��:��TJ��A=ߩ��M<Zİ$Gh#ۨ��W+�܌�c��sh�uW&	�egp��p�֧�zi�� Y�Z'Ϻ�S�L63��}�{J>-sah�b+���٩�j���P� 0v:�RK3W��&+rF�'3! ��Uu�0�@ ~��}���qk�|~ܸl��-(��\\���l!^;HY>�KHkO!�	tǫ��Ѿ��Z��KT&h�R�1�%+k�g��M�]yfd�n&���_�����&�r!/aiY��EC�P�߈}���x��l��L��&���g�VF��_O�����:Ɂ��[�$�#��N6 �̘]�颣���K$�$��<}R����k���L�Dx��;-=��z�{y����7�R�yy� vj�b�|�8?���;�-��o�Hz<ț��ܧ/��U�s+�6�_�]=�oVc�4�U���qI�xO#������, o@��o��������o��F�r)>wACٝ����4����L׷�����f:�����GM�=��w���]���� �E3���[Mk �Rts�����{0�#?�<q����峵� L,1���&w̻�/����e�s���Fu#XK�8t虾
S�f������Z�X�l_�5ԝ���/����{-��":��65ǣb��ܥ�.��
�jCr\Q�`kȏ@m����2���U�dG���e�=o�]ȬP��O��l����^��0HR.˻s�]�j�NGF�g�fxx;�:[5��e�>�&GI<w89g,��!�'�^��J�DK�H�p�<���|Nn��N!?�⟀0��n�#����Xg�Fo�����*J��42Xd���'�&�t��
��9�x�
�_�P.�sj\X��5�;t�#�oٝ_����R'Y���Ҧ�u�,�`��5j��h�}x[6�6���Ak�{�JoU�'��U�8���]l+�[�O��M�u�;M�m��LM��79`7r2;����j|]+8?�d�?S5��]Z�	m����N�MR�㲸��ek�B�N�s����0�H�����Ëv�l�Ħ�%�dL��rf
|p���>��6LKR' �a���"��?z���(�u
L��IA�s��������?c-�C��A#����3���q��^��h�`�`4$��u��{_�,�*�T̔+2�b��S�Mk��mX�"���}.&G:pe���[b;ChB�4on��L'��i��{�,:>�/\��D�X�����~����R�E$��`�QvA̽��eu�c��ޑ�O}�fR�MF����s\��?�<�
�it��(�3L��\WQ똩���f� ��q5: 1�_~�*6��@�1�v2�x��� ˟w(�Iׂݳ��]���:pU�TU����ҧ����J�|�22�� ��֞���F�Ƚ^.86���Ɉ��j:�<�.@b�����syS���s��{�~,��RZ>�������:�,lmMqx%n�=%:a�\@�����(�pԭ�/쐵��T2���4x$t���3%�`����%N��.�˫$�G��(�%�F�� ��;�)��{�m��l(�b?��k�7hC/���-z�HP�(�b��y�݅� ���nj�Pܜ��($R(b)z��Yx�i`5BW�K�-bZ���5�d/��%�pJ�y8>��ҳ�L���b��C��"ݕ�,r��^�j{�p�'��T�n�M�{r'E��>���8���U\�yR�kxs��VնF�\�ԅ�Ĺg�C�j�@c�4�)�/د��Q�=�}q�c��\Zp
�<�S	��|o6�x���$��F�4I�	i���a�����1�s�4p-���
��Ȕ�]
�7C�:��d���z���\���"Y��Hw�K�n����h}˅����� ا`8��ϔ���:^�s�w�������߇4T�ԍ��U�	=֚F���O�t�'2���u��(��I��5�,����xF%����܋'�Oc������ ��	�;�Ó�0l]��-��T��
����]��S-�j
���+J���B���
�B>ipq-h1�	.�X�"E�}�G�]ߡ ���3͖����t��[���X��o,hH����<T��K���K��>1N��^5E��t��Q.�Bb�.�?��~����vD-՗�֍�)Lsmc�(��-��7� �j:��JOI���{mf,V.��V�3�������h%�}$�W�y�2��f@�O�)'��#�oIlaq�g4���r�o0�[F:�r�)��S��aK/7�/��D���R<(��d��pX0W���+�ؖg�d�38�	��Qal�Og�y S�x+m5A��#D��#	]��]A��eR8��Eӈ�Req/�`iXu�QHT��J`Ņ~�.��SRE]oʶYd��_�8j�4*Y��ג�\����{�M
"A���ݟ
�T�U�DP��[���T����:<
"� ,��
��F��b�W�\�T]Sޓ��}��G��xȝ_�e&]B��UjhW�>&H�&ͮh�m�`��n0D�)�A˱ńI���ZO��a��h�DwCϦnNm�#>�/���2�WH4��f��S�Υt.I��,���n@���n��ڲaҲV��aX�XVZ*�G��RTݼ#L�=�@���b�v�s�2�3��ݛK�1��;n �O�bJ�~��DȜ�>��U����h�|�qB�½z�d8�L�63��2�)�Xv-$p2}��B��OZ&��I��e]�<x�"V�bQ\��h�j��l�f���^�<FU��$�z)"y4G]�`n�d���M��~����J�n� �f~o���AD�K�RNEH\�R�N�9�[ls 4b失��Dx?/��[	wQ�-f>� т�R��`�����ۉ�ѐ���l�{4tG��5���X���;�$�ÏX,�Jgܙa��
O�|�H-��z#�ufս�z ��I�5/��HDy���g�Aa��
�}c�$�)L'�7�-N�4�q\{�S�0�/Um.�A�b5����737����1��ղ A�Q�����/9�@8C�؟Α�劘�|3�l��O�wQ��Ȋ�e�-l*a��W����$@�eU���ʞα̷���
Bu����[u������U�P���r�D���բ"X" � '+�jo�4�^��(���\������C��/�6+y3jYq,�o����9�A%;�:GI����/mouyGO ��|Z�;�J���E4�+j��օs�S@�ڒ )��'������4~����F.,��Okŝ翋㙮K�~�q� ���A�6Q]�v�9�y5�ɤ�lM�rY�g�H�ut��$ډ�u�g�*��\�	A��	�	���^W�]瞠x��d�Bs�0�v�z��b�y)i��6DC���l[B5�դ����sXf���}���yᵞ`{�Ѫ��{��$��P����C!�����B���af�ъ`�RQؤh��-� #�.f���棎� D�X-@�+��y����iW�JW�m�(���G�.t�Y�ӏgEbJ��%PB��X�<�?HLY|3��v���[���T���"9����8H�]kG�Y�2����a:r�ak��s�����X=�~���)��=m��ϰ��8�m1����H����j�Ք@7��WL�����������O �:T��|�\�c1��/�&�<ܭ�7���#-]G�wj��ZsN���}���7q9��n����
J�B���N�6�m��u�C��dK-�pJ���g���g�5Y����t�]�}�I�o�j�6�rK�ɣ_-�;�\�4��m���1:,z�*����E!;^����n=�m޾�PU	�Rk�W�2���,�~��x�Z�Vz"[�D)+�4 ����:e���s��7�*���Ƴj��N�i����z*�-9@AV7� �9N�$��c�S�d�?�+k�ֆvSOV�͋��#g��J��TGB��������8�r�τ��,�T�4;ͮz�fƹ����8D�·���<���YS�V��Tp�5����D�|4j���5��ȗE'���\�gh�]�4	-�)��`�%r6�(���Gg��{��N�����p������F"�������f��<�� ��xzWH��:D��Ԁ���I>c>qed������W�]��3�����r���T
�Ի�
͊7nx[���ǳ��9F�&��u"k~�h�ʶ��&�<A�~Q���|ID?9TMZ��:qi���`����9r��3̉2뙵(�AQ��U�����άlO�iV.��A@����RPS$�תvj���]���������!�U[\1���J#�)f}�J����Fv����z��d��fO��}	u��=|H��Sn4B�m�O3��4�N&C��]��d`G��9<����y�i��� ��-�Z1[�����
t�8�|�+j%�`{�����v��\GGC�l;��1����T���t����GCK���%xQ�"��~ڄc1���_O��V��[�Hd��U��i5��˼�����se�<�D�2`�Έp����5."b�����4�l�ៜ]&ܾ9�<�^DiLe��7��$w,ZJ��Y�ɋ��2�;X&�Ise�x��<��"�m0���@��MO�
ʹL���_Té�#{,�����gƲ魉�1��B- ������XWs2ӑby�bs����:���7Q]�[�1@�s<���M���ʹ���'����=��\���-5ث�-�b�[�y��
���K'v:�f��__��"��,*�<'I��y��,\E�)��>�=2s,;��Ď���}ӳ���.g�@�(��0d� �����zH2_`�Iw�������jy����cZ�C�C�[���nQ�6��Djݟ�����ȹo�[�7�ZoY���>~F^S�B��3s�g8��l&��p���p���^0����ѐj�o鮜�>�|L��L/C	HDz���Z|��^0ɚ]�/o���|���Ty�ݮe9!����V��"�఩�m\�x�VW%�f�w�7�: �U%�G����g=�!���b����j0��Bf��&HW�T���^WS�H�����p"�Yi9z���H в`���#c"���宪��-̝�Ή�4����"����&m��~�oyǁ��ؚ��I}f�x�R��o�A��Y�'3��v�}�q����d*nA�L�F,����%fr����=�,>���M��d	�:]�-�9��t����`�9��4���h2.Φoa�M[(&���7�9Y��l08�� *|�R�P)��5XFW�W^���c,��OUI��7t<�]}�2��[w����V���|�W�
��1�վT�i�b ��AdPP��_6#;��+Z��!b�U#e@�=�K���|�q�hR�3CԎũ?��@.�8�@�\�9�ba�}�'��r\h`)���P���N�Ve�2�џ�Ov���c-�qZ�tyǑ���t~ۣӠ����^����!�CF�2}F�|&�v�)�-�M��l[��F�Vm&��E�g�к���.��=����bw}�I���d�q$�9��D㖁Ί�+6%#������g�YuÂ�3��Эס h���ƛ~�n��?��W:�����t�ܐ���K�g�g�������_���6�|ƭ��YP�Α��qMY1"�;�Ir�ʅ~4���R�.�q@��{�&�-��ċwӸ#eL�^�Sဧj�9�F'�aҸ��u�nߍ����h��1M@$Sfey����|fG!����Hk%���>|���߶_���d(aT���GIkB������'/�ٵ�:�sqἾ�@�LSi�=S��g�{��*1y�|�#��4O֢<˪��ˌP	���=m9`7���@�Y�d��W(���0�|�<�>�ʮ�F5�syAX�0��Y0@�S��s͜Ɋ6���
��A��`b���r�����{��� ;����M�m;����n��E�����C;�gcG���D�$�W#{xT�uh K?�v��i��"2��#M�[��F�cѣ�d��Ԓ�7�^��%�q�G(�0��+��\	�|)�n���_̿hu`���_E�8گe��<X�ѓ�N{�-X��N۔1�e+���_S0^ǔF١j����`�$�ZX���;�Efo(0H5L�� тQȆ˗&�<�#mJ`}%4{b�e�Y��� X��dc.!&�F~q�j|9�~���� �M�49m��l�&AZB������s�:Dc,��sr�FS�sr���$<�Ob�=�L3�b#��mIE�>%8H��^�sT��J.�j�g[��p���U������=#/�Pwj��.\BN�j�:�]����	����tŌj�b.N稅n0��h*9���4�(����P������P�#�ي!|��E+��i�0���#>Iz�ŕ�WO?ڈ_I�(4�Ⱥƙ^��'|�F����z�mr�����"�����P�8�������N�.�����e\��B�� x�(W��\�}2�sy k��؜�M��〩�t��a�=�B������'w$75(
)UY���
pE�<�XS����af���ꑇL�n�y�%�Auj������]�-~<�ׂ��l���[��bZ~���z�{�Aj����G��v�kBbX�fcK���)��8�S�	C���3ُ�I��N
@��/�w�L|>��%q��`Т=�7t���5	�Z��r��5<�ʆ@x�ccci�Q��Q�5��_L��AP���
P�Hز�
C���������;���°�6�+����a A���}�g�N1eB�:9H
�#r��O��De�Ӷi����BD�}��5 0V-3��)�A���J�]g+hSg��	nއ:j҈�������������묗���& ��:4h�t��}��t@��0�wȕ��ɔt���E]H1�ogqU8U)��ӿ�:��w�焺��gZ����ΜvŶ�4�/r���!����hϴ�'�%�@�3.�������+�^sYJ���-ݱ�}�?�1]A��)��k�������e�jU�a���P�,:K���$�l��Ꮾ�=8ґej�����DOJ )���i���C��f��������C��R�l� ·�k��"r$�n_��mBF&��b}XU��fG��_��WhQ!{�(�n�Pl��a���xFu5�-��D;]q��jA Ʃ�@xP $D�9��#6�����o����ٮ0���h������h�%����#F�l.>����7������aMfa$�����7+�8�ڴAsP�}�.�|��=�M��*lF�� ~�_ڡ,���HM 2�L-Şv����q���)��n���,h��2��4^��8q����H���Y 	�3�1x����#�F �D�8��B�8�R-����5���d�P��ѵ�����(�N�̘�X'�I�_eyך:TE�%��k���MU	���}��@n�����Xo���>+p���Z�	��ռ���:�>?O!a]�v!%u�}�`�}�t��
ů����$a�+'[׻��am�3h�r�p�4��.�'�hj�l���b"b��b�	�m�'���?ܖ�L"�����L�� ���<y�d���t�.f}�m2�t�dE�JMԮ�4��r��뢻\/����@M�sjQ�W���5�b2���S1u�^`�)�5��K�0r/��т6���~�ET�͕؇6�QyrN�2)Ib���o�Ї�<�C����D�uP�<W�]�8TQ���1���l1ɇ©g�h������}��um�eaK��"T�M��m�LUa�_�g*�=IJ#��2?Q��坉���4]�9��]p<md��h�c;/�u��\;)i8�8A&ٝe�x�s
�f�����E`�҄�חǮ�����'"��!R)>^%�n��1'=��t���oO4�=َ�E�+	\��[�t�m�|��=ED;2n["�~Cf:9p��Y'�T��@����ܼ]��H%Э�Y�h���^�ǒ��}�6����� [� �x���<*���N��ބQ�;G-���(���;�PΧe(��_i؀㍠�K^�6gW.*�HpWbC5�w�궒��ۺCZ֟-�	9#���r�yb~	�c5��ͮ�EN�h+la�7���h��X�Y`</� �اsk����Ս�S�^	����3�z�O��Z��D��R�X�*n����c���2e�r���>��a��\Ґ+�����0�j�����%�T�S���Q��N]v��7�0��}�?���J�����t	�J�Ua��oz8D�)g\�n|�e��[�$v�h�pC���p)%����J��\�a�±��������Zs,FQNc膐&�%n,�f2�;�߽tun�D
P�s��U�l��iBY��t��p��֌d̂ EG��aI��o����8f�G:���g�|��I��x<7��cQ{��Pt1g���l'k�
�ֹ��Ϛ��ȆB
T"Y��F�:ω0�F��5 �Mjt3]�"���7�h�溴���<=m��!��3��e%��.me,�tx�4��?o&�Zo�6^�x����넏�ن5���2�+��9!^�B}H������%N��t:�zy����䛁y!9�:�g!����C�T�5)q�����%�X'X�E΅N�J|�EvJdm�dO�<�������tA�q	���d�ua�����<:o.�D�{pT�+���_�٢�4��z����u��r���|�B� e\L��Ӵ/2f($-�~oG��}+S�ֵ�x�,L���JU�(��h_����IFV��y	�)y=в���p2� T<i��;��]օ�i��~<��k���!Ib�jC��H��l��/���Auz��?��'�ҩc�eիą�bov�� �Z�iF��j���Q(91�2�K���2_��ڭ�a�{�{^c�8�`��2i�>��vT�r�Ы�H���i�Q:�:y��D,���|A	�}}�������frn��@
�Q��Mh��q���j��T\$��4��X�"�$ą���PTk]�z���?d�;F�#��O�h�����@�}�S����C@���C���8U$�hr����[.���$��
�@��1j�d�\|u�薯����CU3Zt�\\���w�	��s9�R0�Y$�@,C
f��Ã�atwDuW"\�-�Gc��_敧�:���WMm��Y���^��؂����ؼ#��?\򒴨b��Ғ�^�&��g$�G����D�t�������:��D�&�^jRY��ZXT�/�F��c���&��g6�"�����0[3K6�52�u���{-A��=#/�
n	&�SzQk7W�n�̙Sر�,����k�#�3��Z,��{���+��2��2��$*�0�
�V�E�o��Q�r/�]���
�N�,�^aI���&8����d.�p����-l����k�1V�Ua�b��c@"!�#��B���$��IX9Yap�
���ۉ��<4 ��Hq{��h�l0M��=����o9_$�Jn �.�!+-4��s.:��.]�"�V�$�p����bC����6D.$i{2��C���e��_H�E�^k��\K�Kz08��u�X|��2_�7��B��yw�h�<�08��|f��N�:T낪�ȳ�*���I������zt��< R�
�^GL�l��W�W\���oh��+ś�;J���}x������m9��$1��mj4p�Y*��x3M`E�Yݗ�/9A}bT\���!h���|)'K�W�gb����U�zL�ݮ]����i��K߄'�$0�4!�c�@cB��9x	�uj�VE��'5��dJ���{qzs�a�8�ˢ%2X�kg�VΤ��Wb3%{���U[(��Z��z��6 7�{8o8�� ��y܍b���IC��'�+�C]A¦��_1�Nӑ]���ǫ%�
s���N�UF2l��{#�+�ު�nc�-B�U��~&�=���D��<�< ��E�:��A��f�ҦS�G�� *�;d�2y�eY'��S�c]'d�2�RG^�Y��,Pe�Y��Y��6�7bY<��7�ѯ�[?�ĺ��'���RGQwS��K�,����j�(a,V�����ء+!�;$�hv-��z��'������5���Y7��"��3�%��]�0�d���n�2���5�T�~�����ʊ���T��oղ�|OP�6Ħ��/� X�]1��9���L�_�+�7**u�P�.��Ӫ�p��'܊�� ����b)&�O�Z��0�?�x�bk�F�q���1��[����}�ܜn���t��sB�:�p�4\$C���K������΀�NS�e�GP�
�pb�jC� }�ˠ�r�R!Y�k{:��>#��NK�H�h��CO��O6b�9�~B$��:<)��#<��H�Bc��C3?]���a!��d_Iw���礁"VcG�8UG	�z�M�����4i��L���^�%��D����B�n�����\��N�0I#^	#�A����#��~�B��4Ǆ3����FK_b��m�3�W�����O�^���k�V�B霰~r��]ŏ�UК@�y]��1Q����}\�Ƣq�X���K.&vY:%ixij��x���:�b�Ï�dK�9�=�t�^
x���m�=�=����Jc̎{9Cla��n� (ۭ����#��vͬg��)aO���$����{=*�?���^ʆj��p`�iM��J5�K-?�����r*G���l� ���@		�b�����h:���uS�'\��MDݐ��gcНG���H�X�V�l�����_��~a�1�}ç�=H��=���k6x��t\�K��7t����/MbBWT��79�޵�����Z�St9����x�o�q�rټ��Q,$)W���q��h^>�� >��okiqT���M�L�R�/���Վ�";��">hw*z��pp fr@o�i8�j��5mhn��/�-�3���.0aL�dQ����CXXߜ�NZt���f�h� D��!>� ����:($e�����3��)Pk��}�o���I��@�ʵ9/a��� V����%�<_���͑���@�o��!_��bD�����49p�pmB��}�{��[�/���p˳t�,��Q��.ܨ�ǁ%�&?���$f@p��@'ak����V�MeA�~JmT�$�wf���GL]v�>��8� ��J�����$�-�җ/{�B^���+<nsË�(.��&-���*8sgݱ��-胝�rQ�(&�V��k��h���6d���D�k{��[w�9��f`��	p�W�!Z�>�)�_w�߲_����m)�mK�aȂ�#�Y��:�g2B]{���/TN��Q&�s�NR�H5�3�|��,�o�u�� �2�q"{�8C{���oW)n8�Umʈ��B�N�+ے�$z��>��M$�	U�jV��L��S��/�� �s���Wm=Ť_�sHq��S1A��{ƎH@�m���hq�]�~l��d �	'���G���� z'�!SaG˙��2��_0g��Y�r�8F����_�mI�>]̈W��B�/�)������ƀ������^/tQQ�3?c�����A]��s5����n��z���iJTE[9�j�=F�Ɲl�#=�[!�'>��Q֞N`Ma�#/��*�Ն�&�����j�D��ֺ�=�/��A8�*p�ۉ��.���,}r��ʒb�|��$HH(pO8���ݓT���n$�k)���.�3��5�Awב7S��H���-�	��z�0�o���8�2��,:�ڛ�h�����E��rݩ�h^ڈB�A1|���#���Bsu����De+����M}���P�6\���Q���n~���f��؟��N�D~�%�wh)�(�.�j�I�+�8�Zc5YN�)Ԓ�Q V��z�Ī��L�'3���p�1G؉�/{��b��]LQe���,_��)#�p4�E�(ԅӘM8/�R�D�'Y	ν,��z��S�����^��\FT�X��y�1S�7q�U�_,lY���aMv"i��_6��]��q�^�ź'@y7(9�7�`2�л�͓�������f_1B�L���dt�,Ou�m`-��'���TFOQ��l<R��O���(�8��K�٥D�q>�v����\	��H��Mk���L�%�D�Y0�w�/r�ͥeV��7
$�����/.���gdYy�Ĕ�������OZ{PB~n~S����V��Գ�U� �z��4f�\�ŕ��h�]`�n����;���Y#���;RJZ�v�},>�.�G�E [�v22�ՆQ%j�Q��~%��q�B�7�G���j>UkJY��J__�D��S�� YW=�������t�����.y���T�@	������:�rU��'��0�Z�1��ƶ
h���}���$PԐ��|�ܪ2�,��	���}�lRS�(Ma<)?'������b偧�Zo�(��f��po�ҝ�c���]���}EHkl���K��&�g�0;Z5�6n�I{SP�D(;��^���;�zU\��d����?x$5M$�4Av��҂A���dvl��I5�D�,��nl���]�z�����g��U8;���K�a�[�3@bU\���@b��A�v��;u۰�3�*����i��Lg�s��M8�A���G�N� ��	8�@k��n�����6'S�rכP�Q�GGVI��&l�%��d\��된��)M���>���e|r�[���f<�]���Av�"gr��K�o�H��|k���;XR�|ϓLr^k\F���!���kR���/�I�Y2�2����![Г��iw�Y%�USP����w@����)n���4�T'p�9)��n��Y+��S�q�*߰ �Bw�j�y5�)��~g��*����*�{�
�N(� ������~J�_H�&��� ���bZRd���R�|/:G��
���LgʾB��'�ڪ���c9����9�1�3񓮒/iA4�C�;�� ��A�z�=��G�|��_q���@u>�27O�P+���.��4�����{�@5�U���a�l�	�M�q�uԐ#�>�Ťr՜-n򌔩����Y�Ό���uPvE5ҫȽ~z.x B�X�'љ�2���i݂��ri�Z� j��;�uve��eW�7)BI����"}I[?�Qa����q,�t�F�IS<<ԢM���4�--�wB����E7\y�"�v�,	��f��JZ������K�v��o?���2c3�H\`�4�ۿ��K�1c��[��с��=����@��K��E=��/�ٔC��.YVNǆ��%�«�>t?H~�N|bqx�&�@L�V�S�`�'Bi��Sk"TN��]�7>HS�)�>}�!*)آ�|";�U���*�g�pU{��5�ʗ���ֵ+��'
�p L]����kF���H�*М�(Ø�,�jՆ�����G�y��71�Ұ�ݳ��X7-@T�1�c���`S�D�W�-��
ه��4��O��N�x�)Le���g��q/��yd�	�Z���B#H����}:!U�p
{�x�jn=����\�Ho�k%ӲP?x*��c1��"����zX�R+VMj,�������Z�P�[�n�9��L�V��*�LM��5}q��!A��Z����o8����S]��JÁ@a�5��K�~ULx�x)�)��t�m����C~)�i/�da��8S+GAZ���H����PO��V�`2D��gZ�n�6�'����L(E>��5��9^����l��W:�|�3�'o5V�9���r�vu' �3|���@��5Q�����{�����S�V.PD��9nk��d�j�(4o���������'��I��P���*�.%6��[�d�L�q0|u��$Y��� L�|/���m�[�I��^[� �ͮ%�-8�=���o2�,K��;��Ug}�j��-;͎���p� ^k���x�9P.9Jĉ����/���U�r@���s�b��܄>Ra�$/��Nѻf R����N�M�.I�sk�55���v�]~�m`�UJ��?�0=��}-tm��p3�7oM���XE�P�`��&[$���P/r�:Ju��T��U[�U��)��Ų5�h5��w")f�ѧ����9��;!��"%����3^*���e��q�����&�6X�G�����zzRN��D��&������W�/�q 
��1yr�F�"�Ev��Y夕+N!BǑb��2M��� d���
|������>m�άhRw����s�[.�b�+D�8���u,��^�^cHB�pl�!�.�}����9�D:��'Ց�
�65l_���@3��,�+fG~
iI�a�s�B����̶&^�:l/|6n��s��P6��Z!��D��2��#R�z4!���o��'�j=o�	g��,ZYz���	G���}�`�X*np��ؾ��ݷ���cR����,��-�cQ��.,*:�'&��b�%���3sԶ�M�4�s�r��Y��i��"�y���H�E�P�a���8��܉���%�JA���O�lT%�p��1VlM!�ʊ�4�t�lX��P���n�vprk�;�Q���5�Fǌ�1U
�ZS����A�꿮�6��^�;T����/�Ÿ̏�[-X'06	��& Ț��P 8/x�/���q�U�,�b��"	��#R�X9I�V�9Ȏ^�z�x7����>�J͟�4Ix����b�^�6k2W+�o�"��R�:�Lr���!������}�xQJ�W�/�{9��<X�x��Z�8JR��16hQ2B3u���G��f�?ݜ�*0�����-�0X�j+S�������y�V�~n*�&�u��n������n��Pj�-�()E`��z�E�-�Pf堌ͼ&4�*� U�ݰ�W�.�3FZ������ϫ��VJ��C�jH�ۻMٽ��&S�w�S� �����K����jP\�q����d����oY�BC����A
3&��PYr3o�<�	 Z.�9�9V�
��?�SC�Gj�W��h?��*=����J��a4�g�5&��g�fc0�L���V<p�P�.:L�������H��jz��z	�0+KǦ�Ɇ����&a�]B�8W�8��e=�^67��G3,�:a���$sė���`��!�<O˗x�G\�a����u�o�X�J־���fv��QV(�:G����A�-�B����NƭŴ�&���K��R�B}���P�i�� ���-�0���!������x�Hj��d���\�U�c��= �]�-��VmUCg�:@��8�>.��4��������R��.���;RN7J���,�v�C�<�� ��@>��atd��r�m�^�[8�Dzf(�k�ͧE�ߡ���_'�I�ji��>��B̪��lҥ� �i�'=��d��r����N����[%C
Dv�?M3�ӄE� �2#��4�2e��;A�(�%1A�A����h�6�=�w�ና�D|��zV�J"��`&�g�1U�I�'��!z�ԛ�7���Vf�cYe�R\�w`�Bz��+���m*H��o4�����E�U�!�K�n)œϪ.���tlv�(z%���>@f�)����/�B.g|s��X�L(��4�>?y�kH��l8�z��B�L}f(+Qs ��^��+�10�DǊ�<&B����Y1�=pGA��ho���?,����]��ȓK8���W(�w�=[�0���~�b�2��ުO����x�Ń�s��p#*!mj �pJwt��$�lC�!h��]��
��Jz�W֎N���+<GW�
�bZ��ӕ���\ؾ�=F=�zrfy�y�4����f&;�n.��3�p�3�|ͫ�"�(^��-���b��֮�P�*w��D�Sn��)7P�d�Pu��p�ź��C'���nz�L{JX�L��6��i
♟|E^D�	�B���8�G�I6i	9H�oL-�ᰂ��E��F�r�,���#��]�!���W�]�D-�e�����c���u?F?�{��Aם�5-ey���AՈ��;q����Z=G�H���LZ�N��Q٦{l<k�͙e@,jS�ZS�95~�8H����GЛ1���U2�W;l YkY����,:�+��	!f�⇴9ⰣH�6��i�Yk���滃��S��� o+��I�H(މ՞rJ���Y�lt倖⛂#N���]v7��S�����(��8)��olX�E�@I3B��>Ї��\���:_�^�C5c+�z�unl��Ǧ�MG��\�j^E*L���`b���'�A��3��6C���[��>s�Y7_�����5��<�#ʮ���I��������x.�� ~��.�l��R���!�����m��G����t6���ɵW*d� ��R�X�<�ƥ"Pց���9��G������?�+k@�����4�ŕ%�g���;9M�כo
F�l�@�弃���{��a�0q����0=c�Ȍ{��6K�l�~}��s�J�CK��=��e@3}�,�̾#�SX��荬B���R9M(VI׈�-��4�Ub{d����V8��-Ur���.T�$���7�!"��N�j�Z|��U!}�Ur4ļ�+:J��5��yK�o�wo��e�7�m�s����&U���Hq�Pn��.��H�t��7���צ��\�U��%�)E:�r�����p�N�Ȓƾ�B��c����	���<���$fa:�~��� �r&Bi j��RsL�Z8����{,�#�~�E�Q4Z��T4��u��=H���P�,��c@o赛N��]Ј�[7X�T;ժ`���lG��hi�?wX`�R���s�'ϸc�Z��EoƧ���۫�`���ؒ����Ӵ�Ћ[��v2M�%ʩ�C&ޝ��;g�`K�;u�$����p?el$�}��XEZCn���`:��n�>�2�|!�C�w�:h\�3͂�Dc�O�][Ѳ�����j��k�f��"�j�>_5D�~��lPぁ�����FY���6�������b
��tD��W��M��>�Qe9,�lv1�wѽc>�G�������覛�X&u����i��&V�Z)���lxW|CPV6�j�@�W�׈c~;%|?�'!T�Q[��/K��x�q��3V��_��^7ڄ�b|�V��a��"`������x�V"5�"푊�A9Wu�1!p���&�����He����۽"�u�	+UZҼ�Y[�c斠�XPW�^_F	�����N���A=:��|�L�e�6��㟛EO=�Y�4���Z�g%������L���o�=D	�œ(�D��S2��1����8s�p����%I�~<2J�D�
+��<R>w)Q�ŏQ�X�r�#&$�ŵME�j�=�0�z(,�Hm �)9b��	�3S@Ƞ<���6��AP��5u.d����@6�N�sr[�\_�ă���9��?;
lb3�q���1v&��*���2F��oaU�$�7���H/�������������w��Fxkq�R��,���ZI����q/^���/�O�K�T��3Mcm}�U��DƱ��C�����ɂqL
�m��JX�7[M���NL��	r�uL��J��Pg4�.�/�ۂ���-�߆���k��̎���"���N�d �p���ځ2�	��)�CUĺ�p�/�U�4L�Յ��Lpw&�ܯ�ЊI��F蒟3I���U~�������<>v�R-!0ﻪ<jQ�if���y��(�oR��y~e��272�+�"�f���k�'C����L/]3�^�C
��D�9%�9��ZKp_���(H��K�%+���(���H���[�,J�;�voY�p����e��I�1B��V�b���'����i6T8䃔O)�`_��q��<&���kV���;p�� L#<n64�p+�)��B�D]tq���ŝ�U��ODI���RP��A���\�GF��:�5��ޙ{S�ٲ��<�C���/튐w�֠����LY�M&h��b�mL� ����|��Ix��sIJ "��i�F$s�,�sJc��HZ�ѝ�h����&2��mI�A��|��-�mUCj�*U�/�S�2ǫ��~���ۭ��u�c�]?��|�R��7�N�Sӝ�ܙ���q�d��9-���Ar�C�{�+)*�b��	��~(�ʑt��:�E���\���q�/��;�H�q�vJ�VP�Vs*����9W<�����P(2��8gfQw��G�И��i�&7��!���ŌPFJ�c�/}"��~��!�	H�9?	ԊjiW��ځ�E8��"�Q?z��a���5��&RH�_\�8FXn9w_�����\A&���� �m�f�Z'��aD��6������r�K�����Z��J�H�bE���(��c�do�r� y ����q�s�VX�A��<>]�x?��~	K�c�8E�b���m��l,?{�b�2��wT
cl���IH:ĎC?�wLNέ�:�@]V7�G��=R�V��#�!��NMK!�����?�� 9����2�e��+��R�qAN��e��*��<Q�]Up#��a������H�k�>�X����<H.w��g%|iND�vqP���P���ǖm�O���2��os{����(Ng	�w�u+U�.�a��WmB�4�P��aY �)�\��W1�,�UBa��<L����&��f�j9�d.'������x�m�=�#W8��d��g6���T�/����Ɠ���w�'w��+���]O�:�&1��b*�gI��ԗ���Ͻ[�#\*vow��1N�o�=�u$�"�mgV7�)��'�,^F�
�I�ժdj�' �ˆЕ��FFeOߜG-v8����&���.T�c���N;Nl΋�eYy����\��OO1���������"�3�������#"�3����߹������znt�8�ދ���Y�*�ե�,�u����d�8���h�,Y=�i@@v�/���z�4V<��U�b��i�}A�[�`m���^���U*6�ƫuJ��\���f5�T��+jVŶz�����[ථ�K�gi���;�r�B���`XS��!K�hCжzr޴��@���š��7�U9�sYB�hs�L1VF�MM�VM������j����`��%�fy��.�PFT}鶅�吡�L)����,�創Iw��ƍ�<|��S�6)�d:U�癆�k����cҥD��AVO�H�8i88*'i���ͤd�Ǳ�sl�Su\�q"Zr|�E/@�)XH��?�4w�tzM%�����	�_����۰�_,%��~��*65TQ�ny�a����q+�={�1�۝!^R�l��@��|��;\���I�� ����>��NW��~sBOm�^~e��+/u��5ܲ��ώ�q���M�cA�NS�$��WX��ZB��aT�cUK�>?���k'{�|��%�M�ԟ�Q�eI�.�W�#x�;�S��+r0�T[I��Jb�}o#������"| ,�.괼���n��"6jaKƂ���ZC��S"G�{�2z��I�g4���	}�櫢)S�|�|bʬ��D��t�����[�nn�P��X�56��P���Y�-�Y���[,TQ}�c,�CO��`�n ��c�ી��S���1�a�6�\^�*�W�म���>�<U����3"�~(
?��1�y����/�tkcr���1��ֻJ*�X�$_�@��z�� [��V����7VqcF�(�7i�L�dyO&{PVXYM��A���0T/:B-:T�Y�H�X�8�Z��(��ָ����KCDfI�՘��h��0Y��8��p������@
�!DK�5_��Y��~\��{�6�v�'�]�Z��Rr�U�S��$U=�&�Ffȑ�5�I�:��.3�l�4s��6+)��8X��;���ܤp<J�G	��A�U�0�Ǆ$w���5����>g�C��~p�r���t��l%��1΁�7h7!��y�A�
0!F]�G��!XdT�7��L��um��B�ߤߤ?Pआ�R��R���Ξ��!�|��=�4~|��'��m��R�WgF���krF��������Fu�4s´�Z��G�l�쨱�F|N[����a���㷎��e5i8��^��%�	���@��k���=�0�fFY���br\5�H��m������fǬ���e�L��Hܐ'�)
~���W��G��f�K��mp���c���#�;ۉxx���T�o����TT�)�����Y��z�a6QV=۔w��8t��K-f���/��~�3?��s��oz;,���4���o�5�n�EE̶�3�0�@_; ��sȽ�5�coy�*�t�4���5u�P�S77��o7f%�?3�qܦ*'����Y�oy�|��2��������P{m�uȖ�}��T�SvIA{�!��zx��,��25����ð8m�t�1�Y�X�����Z�d�y�J�� Yl,j`������}�����x$ ���ovYY��]+q��HP�u�9�?�pg�Y��l`ס�W�9�ڦr�����+�ڡD�����$�Ƀվq+/�d� j�Hh���)�a�o&n4m�jJ��N�ϫ<�cR��!��tD�n�8�O
ꬭ���2?�wV�F��
�Z-A���N���]  sA�#�ݾ�)P/�:���M�+�� v�����l�~6~r!y�3�ʊY��ǂ�CR���,tX�Թ�W��hl9� ���x`눿9�!�{"�G�2�;3䒤$��ǰ6�lF�l����FN~�y���N$])�A4�ձ KQ��`?�HJRB�{�G���rPr��M4�ҌW�*-�+�L�S�-�-��$	���#�ǲ��
�<��-h���c-��ݘ�q��-a(��<.�
�����i��}d@k؜�
�S�Ƌ0r�7�ev4^�/��3��>���鿳ӯ����o��C�̱_��$�!�&�Zo��*@�o�j�TS)M�X��̵�fӆN9(�1�͑i����iq]�7y�h?�E՘�w��(ͧi��g]Y}�tT�P/	��V�ح�7 ߉�KJ�?pq�>�X:�,m]l{��@�sP�{�+;��x$[Ř�I��A�\� ��o]QL���:p�S��}�vc�z����.
4p�)�5VG����c�f��3�7���}��e�,�K'�v�)�>m����� 5}���p4��2��t��B�+����[6�B�~s=re��5������e��|�L���C���:�]��Q��}Z����~�Ocr#�UD?¸!Q4�;�l�PVD�"�9���i� v���p�dɽ�C��i4�L�X�w�5��
{��9���U<�9���<��؆��v����g�P�l�o�ε�`�-)T�|���`�Gmn�&
��/�����}�32�VgZ�_�L��"2����� ��k�<K�ἧ�γz~��?Hܻ�0m����Tc0T4p]�1R��~�6�G/`����d��IO樚A	�#쐈��P����\�]Gп��{��I?�9a�$��(����V������B�f
PF��^/�b!��`��ĩQ�������������U�"v�'�Q��[�gƵ��	�y�v]縎!�����{�p׷�C�	���i="��r+ӽVC�+l"w��ko�n�� 31'P����C��Fy!�'�b�uۦ���U������F/�3ZX�����i�41����z���(��edY]�k�	j,�M�Y�.�9$�g����cΠ�]$��lq���A�c5��*|��cd���A���yc�|+�u�B��f�)�n��̸T�q��+�E�lC�����#���>_�������#8[���WK�=��a�Һ�i�`���WJ��{{i������[�v��/2��~��� �
حNQ:�j��R��n��N�S�8#��{���k@7X: �=��$�vmMQ�,as�mm�%�r�)��ݐ98G���ASr/�k�ذ%�[�M��m�k�#��fT��O:<�H G��(�������ɑ!�k�x� _
͏�D.�� Mc᧔%RUD�|�2�~)-�������;�w�-H�h�*���e�xn����[9����}�(@�����N���%K8�V����t0�Ƶ/�n�I�s_��Q���tio	EPR�w��"oR3��S7�l�>�U�H����<��A�wdl�_ʜ���Ң8���+M�8,j�9�kʿ�?/�+��ʊ��4��e��������3��q�[����*܁��LO	��p�r�� _��m�z����/�Al��G�g3n��KYU��Zl vJ���&�br�=�W����#��:�8G�l�1:=��o`tYA^1�p�OSwD��:%ZR����?!��m�bh8c�~�=�}ք��6يP5tF�l��ʩ��ۻ���tǊ+<È��uk"��Ǩ�װܲ[�l^In�k��9<����k������a���q�Q�4Vgw�D���+ydR�h[eɐ�ӓ&��ģ�TD̮��g���A�Ĉ�l�מ�u�ǃ����@�#�O'S �b�F1�Dh��s�}K$
�P��9�	f#�]r�T�@e��f(8���'�g�i�ZY�A	��#��BEA�wC�vy*��]QZ2�
�� ��	գ=�������xE�l �K�;�]�*}�C���Ib�e����Q��	Z�[��^�З*9]ډ����`m��l�Ht�]���m�m�)�a��-�/����i�ncP����}Ѿ}���/.�
�Ңo=Ԓ➇G��K�ȓ�ɞ:dD�\�(���.I#���|�ECֳ&�M�����Ӓ0ˤ��� ,+�}�+�ݚ���V�p��8B�[�];]d3��V%nޢ`w�#cۛs���eZQ����YD*�ѩ�?Fbkŉ�.j�����_M���k<��Q������JS&0��m���\E���`B��<���1?��3
>E���h�E�_��,}:��g���R�ZQ�]ѽ4�\��(Χʩ��ڿ�>���A� ��������"��	���-s�`�n�	�h����̔�u8.Zj�Wg��cBm��U1Hx!�B^4�ie[�O�nK�_V��R�j)	A��AwF��HZ��j��B�̕�����竃a��O9)Q�\��/w��P�B@#�jZ�kWGL
��Ŋ������14e���DK�:L�W����;;���U�%��/SH��8���6�+mzI���Hh��k�xK� ��K���, �'Mx�����K!S�KeC_�8�\��<��w���7���܀ChR·�5�$�KLw��m��#�6�.KZ��'2����I;Lj�C4'a�E=�x��}z8��M<��g%*�n��]ͧ�k��&|��Hr#H������h�o}9�Ј�y��|�M�[�\��j�_��i,Ž:XT����^���qB��@Z�:C9��$Puzte���L�O��d��<��p�ǈB�+���b�%��aNrB�a"&���m�s��ut�Q�͘��9����aH0O4*�á�W�r�_����1z�����!�:�4M����̑��;��~��,93e�j�Xp��t���	6'I`-�g\:�m���a�U#��F��~f0'V!���6}q؉wO$F%M���y~�|��*"QȻ�F/�=�Pd� ��V�$:"�2��|�9�KPHS���R$�~s�`1ф�v�D��v�
� 1�S�(�l=~��6���I��e� ��GZ�IbCĸ�˻�%\bu�V�5������Ԓq�ySL�B"��^k�\6�/�j� �ߙ�M�]=R���g�C8���Q���m���"]!��O�w�@�2)ux���2�Kx>HQ�onث�(q�sz�E��c� ��[:8n~E/��|��7�_6�R�,	��#)R���A��̎	'l#C伞\� �*��"5f�X*�伄�{��?f��� |u�a��/W�Ă�e	Q��Ȏ�Y�ˬ���␲)g�:8h�����1gY r�����Vк��f��T2{f��С���mmoeg�j\�P Y�TacdB\������ps��%����s��z&�r���.��S�b=DKg�&U*��ύu�10Tb5�+�1
���>q��ś��آ�^~�k���e�]��,�C��)��1+l�%�l!O�fu1�[$�=��\���"���q�����QI`���Lwi���OW���E"�B�~X����8���?�+�2����V�%7��n����r>�v�?�ԁL�WwPE8fqS�Ղ�7\,�^p�����w���viܰIr�!�M|�k
(��R���%�?�Ӿʢ�+��q�W��J�0�IY����Jeسؽ/���S������t�0����(]t����E=�k�NIc0�l��uA�@_=��)�)�C���#�Չ�{��3��_~Q	!H�'��b�#�I�u�ڑV�":��Y9Ѷ�����L>�T!�%�;]*��<�_$an�{(�cer}<2śq���cX�x&�.��{��V��i�"�.$��KY۱��S�d/����?��o!W�H;Z�1Kjא�U�L�	�G`ю{Qs�<��pk�I��-��k"�%��[`���=n�XD�ϠѺ�{A�v�����������*��B �{��ТyBF͵�X�Ut(#`�6va��B����Dl�7~	z��7�@Vt�0&ۦ�ӄ�X�1���Ȝ������ŝ��6i	�Т	x-�#e)	@���R�?��>�tl���)OۓtWdZ^�
������ A"����l�Ԫ�o� ���%w��ibZ�h���݅�d�e����IPθ���j!��!^ו)�������n�-#���鐄���\�`H%��-�w���?`�G/r����C����Y(ĉ"��?�OѸɷiE��eLA3�_�B��{���F���C`F�A:l���DςI ĥ�ʽ�l�ȗg���a�D��l-�Z�y5G��c��K7W�#�u��9фV��}��y6���rQ�~�)��;5���E�e��׀|;�h����,�Ն�= G�nI�|�aG���+z9g�)cW�US��h/{T@"�`�zW�f��E�����w��\�o>@�Q�m��6��׌�&-y+�r����=��J�x����^j�6�*��f��!�(�Ti���	|UP�µ";�L�q*����o�e�>_�N��j[r�%�^��܂(�oʉ6�*�mM���8I�c�'�])�����m�l�Wؼ@]W�����[��4���g����'O������)ģJ�d�if]b��V�1K��j��hd�[r=�#�
�L��b	�%�fM�e��o��e��j8�}l%�&�����˂�G�2��b�.\$b󾢩0	�-#���fJu�LzDXk~��+-,��q��f��'����|2�&��Q|�o�\�	;?j�$a�Z-]^��ժG!�An��ZI�e�u��+��T{XR���!��̃'������2�c�F!l��ˤ�C���+�'S/�s��F�i+�����VlW�q��˱t�.��%�#хa��QJ�N�����$�J�FђL�!}W��!�`���V;zä[6�'Yڃ��{��������&OK�4������t8��>�5�j�-Gk���J=uw�mI�(�2T�-s#?h�;=j��H�B���m��S�?<�4b����U������9���x��D<)����s+M� ��8KM���秈X�i��~9aܵ�a�Dr��h}��E�o�M��f�66>�%�TwYÝl���.r�#"u.h�B��<��o�j�'�%䥓@�^�<S���F��i���r�cyI~!�X�S�̚I����N��F�-���S3���@�vWE���Pv/Q�`��a�d�/|8���K����Oh�$l���6h&�>��M�sF3_��io�J=��}��A�L��L8N���?��x�&�V���^/H�!B���yeB%�J]���Ҕ=��|JP��Bk�]��J.��l�t-Nz�}:U���L��������z�X���Z�~m�J��?7�U�c�w }:���uP�T�+C�5��l�� 7=��,���� ȝ�yL���eM q��F�Zx��>Y���=x^n���J�5qI����`�7m�/�X�=aϷ�#���,Cӿ�쌲3p/�� ]!�g��xɛ��]�%s���;���k��+���;�xee���zd��|��TC'�cƝ��2�-��Ԣ攳Rt˓�4�5�Zp/�},l���Б����E�����U�c�_�T���?�!!{|�D���i%X�a�㳋_����]K?�C
P;�˴�ѯBs��� ��9�b�EZ���?NzZ-m?��c(�UҜiM��2�	3GJm�B=C��`��o b��D�"��EY��k���/~J`��i�L hޕ�<JY���X��sy�g�����5l���}yF`�|a��C0���D��X��s���a��|����%ʪ|���q��v��χ���:�����n�����N�~��,g�Ҥ���8��nSc?2�6s��ʬ�(�����Kp�D�ӻ֟�J �~�)��c^N+��մpW/��ϑ-�R���ꤹ#���sޥ8%�\�=�H�f������df�Ȱw'x����X��"�,O�K���b��k?uG�EB�����v�ן��݅��Dٔ�'$!��b�7Z]�y�I{@��h��K����vċpj�M �e>*���+�d���(�O�u5��E][_��4�Y/	���A���rؼ��F��Ƽx��O��+�����l�EPX�d0��(�P�BU�e�*�)w߷��6���un�L8ݒ�22�)cP�Hj�������:|�f��Kͳ�U!]��%ș���:�Gw>����F:��K��;�.�����|L���rN���\�F��m���3�Q[��_̟=_��C#+q�-��n	��=�=�8葾ʰ`�=�z���R�_�����A$�i�n
8�Y���Ʉ	D���W�# H�ӔUJ#6�[S��ʈ�w�Cg�j���3WY�V���@�s�����-S���G�C�e��/:?+�-㯈���t�1��Y(�ﵴ��� t�÷^���g�fF�yC��>`1�[���ބW鹟x�}�����;�J���M7j�?~e��%,������-�ӐǌR�T���=����\4������Vom��������{��-g���&Y<C��	�Q�ً,>^_!3�)�k��B���b��S��hTz�&1�-E�ܩH���|zNa�a�HҩiGwD@qm��Tc�L�X���H;�8�B-��F(kd��1N�`[����_�[���4�\�;���ppA������|���������=Z^f�jEc��~~t>m�Zr4�_aq=����
2W1,�B%L���m6�勔RTb��� J�oj�BU'���s�+䰣��cM�\�8���紳���W?ڹ^Yy�b�ޔp��=ZF����ŵK\��ַV=l�s�V�Wאw�U��U䣺��9ʍ��f��=��\���J��䉇'i֋����#�]S�=r���u��.<Y�@�W"�_`w��T�^XB����a� _�K�:B���>�0��x����6��w����E��-nk�|Fհ��p�'NV��w
5�2�����J3�av�S-*�U�?�q���#e_+�<5g^�RM)�6y����0��yh�p3����B�D��"��X�� '�}�.*�P2:�(��/���5��F���=^��������w=.�%f�!"�ˉ�v+���Wa���l�W�F�P���+����>�E ���Z}������|o0�Ã)�ZS����O������c�fs���]�@ �]�o����'|ft�!�JLm�Ð�PX@�Q��e]�~���9VSE���=�|�uK�쪿�DD3��cT(�����0�a"��37U1D/<��&Q�v:�;��-�
�ʭ஡������=��=���~P6�m d�>�6%��^ͷ��f-+qf����u���-^
eM�.� eh�qf�٩my��<=``g�?
���/���B�{Õ���@6C���gE���ڿ*aM����0��6�pYN�Ͱw�=����\���u� 0? -���^>-�+W��o�D	�!��܋A�F���x�r���I�ا��	�q���o���U|̬�<�dQFL��^ƿ�p��&r���X^^�5eP2���/�^LR#�<��Zߺ�6O�(?�?�|�R���.��vN-��]��W���72p���	���l�������8��ځ6]�� 0x�4���f�������T���c[�E���M���!�)��&i�4���j�αИ"���o�A~��X���q�M��O��G����8��G;N�!��6ő���ѭf�kljO����]�%M�^�l�;�1�&��D�t�`��e��i��>��ԚhX)�V��~��BA����r�|if˗�Lr_����X���F\7p�g4��1�d��CS���J��uH����N���I�4c�[Ь*)7��y��1�jY�}�0�='?�"�T@@�4��Ps m���{�\�xi�Jd�e���7��z�;��:�UWM�{*��5$1Z$��DB�3�l\OU6E��=�Y�N�11|���A��p[���(�����8ӵ	j������w��'!?L��`�$��xVP�	������7.>y�i"���i�߼^�pv�ou�H�\�
��p(%���ב1�	�u�[���`nd����X�r�WKd��w;�q�:��n3k��݆�*�����b ,�W-l�iZ .��3�,�/�1�c��.(��̌nC�ce��	�n;,��ˊ5�����F�"�_�l� �ix?g�=�!S�����.�ˬ!�E����c|�ጞʸ�7�2�):��3_��Z)�[�{��>��_2s�d�"Br�[ ;,.:C�uS�����1���Zd1�[��lk���x��B���������B�&KŤ��G�M����E�uV��_��h�w]�d?�8�R�cv!��/y�����>��zh�㰳;�5������,C,��ɚwA�@��4��<�#,1���:����y���ga//e�m0٩���ͱ}(��@����R4/�A!Y��[��y$}�>��")�Bt9Ho�P��7�|��A�ښ	R,�������ǗRuQ�D��=�	9�W}�ԫm���������q�#Vo��B8�~L��J߈��6�"2!^(��n���@�(����T�)�Eˏ�����L����H`��<�_�l����d1Sm��ÛG��qM+l�f� �J ^*U�vZ�x��z�S�.�N�W��&X�Z;a���gک��������M�w�F����R�_��w��ո)��hD.X��Ȁ�g��I̫>=p/g�9����?�0*�{�mR��92��v�;?�qͫ��~* [(*M�"��#kf�v�~7�g�v^�mfV���m���ʛ��!�3�8g����R�=���i˧�@�K��'�C���x�r�A��ÙuZ�I���X�
��>C�`r� �~<�'��~��c5�Pdu�ְ��)���[��/e�zX��r��fm$��kΞ�kHI����+c�A�^��q$�v��4���E�xvY�h��K݄8�:5	��'PyQ��3T�k��!���K�t��3��F7��ٚ���ax����r����x�̒Լ �a������e���}��X+��%���1r`3�^�	����A^����F��m�u<n��C�*�#�Ŀ��n>�}"xǕ�m���"�6'|d�N�k=V|� �����{b�w>X���G�ܙl�uU�1T�j�Ěg���D$���dS����O���m�Lx�,oXf�Ԧںk���΄�U�rk/xG.}��������Ra@�����ˍQQ>�d��9寺���	��y=��w��w�j�v�x�}ܜ[�Q��&Y	�y�Z�y�o�r,Ɣ^�4V�x���}I3w(h��b�>xs�����_>
�;����	o��~��2�%�!TV����c���wc��W���E�t�n.��f^j[#Ѿ	(����9A����sJwO2>���tG_����E5�V��d���X�s���vѝ�CNw'�m#*�+Q���̒B��X*{�����FB-o�S�� Ϡz��*C0�E�n��(l1���?3IZV�r��P���{T��D��1Aqhv&:�jo@yRTk���E���.,Γ������������Ԁ��*�E>�u����׾*��P�$���=m�*��xp�4$ A��p
C8r��P�%rp}�����$gˍ�z�F9��|w;ص��!�+ޱP�r�?-c�D��C�0_Çjݗh��n0q
ھ�� ~�4�=��L�MAH�i�2d�\���v�b�>x��G&������R;���z��#��L���-Z'��IG��e�:CjVm��v�J˩��ITWේyD^%�7�u��S���{��{�ž�ْ5z�]���Q��h��@Oe��n.4�0\ 4$��+����깄KXu�bM�����2B�{c/��{ n� F4+�Jy���H���?��/��C���H��w`9�5Z0Y��&	4��eku���h����#����X�0�-��S��Ƣ���X�����]�K�E��H�s\)P��2/�z굔b��?}h֘S6W�x@%��|�6�����`�C�������CXc�Ej�����)��
��+����C�
&������I������_�7�K��ʫ���$����Jh�*��T���p�$�bUj+��oB"kKb���=�
Z��`רĘ
���+���t�'����*�≫�l\ᱜ���!Ȓ�t��)�)j��{cW�(����9�Wy�\���U��lGE����t�'+�����<G�>Qie�'��l��<y��aOi��t�X���ۖ��&�8<�_�R�rW��Q��z�*gy@�i@�sC��$�?� ������\2Ũ�P�>�h��`ᰭ�ӌ��c�|�+�ec �6��א��V�uRZ�/��C�9�w�=���8�W�_�
��ot4��|+z
�p��%�����,�*h�p@����J���K�E�6K��$�q��Y &��
����(q}K�Xk�"�*�#E����sl��Fv܋��YN-Z���U��E�.��yN�i�O�����8C]��6_�`x`	\�3X��OL��ʧ�{��񹙗���&H+Xq�يΟ\$��>�#�3>?�&*�-�c���r���Gwy��L�x-��Dw �q"p[������%�P��<T-�
E���۟s����،�#u�~��O����FL��rV���9t��J
��4jθt���MC*���:~����?9�|�����ψCxr>���v�j��8
�=�xDdʏ��8�����󖙍��P-~��~Df�N�/�g��ӛ;!���?��n��8ԣU��'��߭��]�d�q������`��t}��.I)@�O�R�Ҳd��1�e����'q�5�n�h�zͼ���:��,�KdZq�k(�K� "X4��x�2ธsCo�9�]	`R�K��PP2���TuT]�^K�)�e�R�	\�8x�h�K��g�?C�l\�K\����ϑ��KH�G���)"���z�x��j�8&5��*H�E6�eN��fx��n��:oہ���shC0�%���Z�'.���E�K�;�?�^5f$�)A2��mAR�E7���@�i��xn�2�QU�_s}�J��q-h��`�������g����7F+����i�Jr@n�Y�)􇲱��XB�F��V��Lg�'���\\�-�W9�1���oC��gV�t����/�=|�����UA��+�4ɿ^��5�50��M63������:XT*�*y����c4�����g@o���7����g9
�ϛ���kS�n���k=?��%
5�I���&�e�..��n��B��������2�hL��C2����k��NBEe��^���ǣ��9(�#��@�_��!	��	�S��t`�=��>��%q�]�ͻ�!��f[�����h����A�
�j��&`t$`��j�?Lsll(�� An�վG��R�$��q�[����d���
[���K��;o�<��u1�5HEc!�[;��>���&��]� �m��z����ҙ���$��D��?@:�'�c����V�ce9$/:��'Te���M���UǴ����z�OU�&��ɐ�F�d%��1?/� �>�t���.�|���\�C���Ų�{�]lL�b�%`o��m���p��m��N\ ��&����h�̻�X�*�� ��zԼ��N�j�|��a/4������S?���|��f�L�7h|�i�r�2Ot�v<QB�nI�x����}� �7UU�tox����T2r1�w� ������I�t
t>c��q���~_�eS���J�p�M�V�O�2c��cz��1k 7\.��]�Al��# �	��K1�aZQB����Dlv��P�����|�'��Qr�qன=e[��(<C�ьn�n��3P\;HE]�A���/>R9�&4m�0���|�H��qS�̫�E\��6�EyEX���PM�������^�ѧp�����	4R�uō�%�k�k��Tg���9�[d6�x��|ރ��K[�L�\��,�wBJO��>	]v������N��v�x{�O0�O���y͗U�v��>���pͨbY��GM��P�@�W��=,�{�x�N�X�	���mm����(����3��܀= ��r^W��`lb���6���_G���/غ���3����Ѣ "�Z2�s�v��`�V?��`dzv�
^5�E�a�.�t�%�vmn B��%��f8���	G�/A�����x�~ݖ�r��U��IA7A2�%$����uO���H���D���)�0@,��c�,�
C���Ʌ)��+�:��e�(Ec��ʪ,��mA��5W©2is��I� Zɯ���`v���쭊N0�w��ɯU����&�x�ݴ����q��O~�C��g��q��CCe(�\k_�r�Ո�]���T.h� �n�+��U�K�r�k\�C�ʗt�]�؆�,Xl�ϻ{u3��3A��j���C k4FDrw�<���G)7ÉĺL�Of�2Y�4Vrs����w��o�͐n5v8q�-�y�+���Qܑ�8� �`=�س��I0!b&�{,����'�*>�:TP�	��h�&#q�����I�����'���Bo�	�ύN�z�B(�~��ʛx�l�k�[�M�����.83Ԫ�-�O
���x��߽��6x�Y�InⵉM.j5��<IB�����(|~�I"��3ű�q����$��w�U���a�vyx�f|����h�q�1R(��L���_i�^>Z�b�Dz �N/��>���eF�Eeڭ��:!��H�Դ@��/6�dL��90#`�G��j#���W���r��(�>)8W?L���X����:��b�h��u=�Ǭ�ֺ=wo�#+�Q8��kcQ�ig����y�v0���u��:�+�
.���f�q��B����T�#� ��:
�/�*m���!�S�O����Phh���ھvʕ���~���__�P�
�ȍ
xW���8>	�>j3j��X�6��F�̣M:<;�9�D5�V�h���q�X�_V�@�lK6����<���L��7��*:���o0�(K0�h�S%�"�m��,X�%���;���8��j@���Gֳ�E:i�y��2�E�DZ����,���I~ʁ���<AG�	_�\՘ ��Cl1c�=�*$j�E�mA�4�Q@��s D����>)�C]��Im*K�OYd�b�X�C��20Dlk�/��F�e�;���k�D�)3�jyT,fA�!�vp���Kя�)�^\L�au��;�=ު�ۜZ���Q���fz��W_������u5y�?8h������<��9�'"��y (�Uw7}q�&+���S�~HE�DJ�pz��:��RG̈́��P��97t��m)J_MdY՝n4�Z����<����|���]!O$�2F��ۯ-���Y�N��+/
���AX �A �uQ�h��fn�4���.J������3(+s��o�G�"�t�uƞ�yh������$��A����!p��2/<�o<������Xm�Q �lܝ!�ǽb�����c�y�:��F_<{�/FC��,*J�֏@�%�̼Ҿi��g+L��gӅ�j�GB�)�ah5a��e�3j�e?F˓N�����p3�t&Vhe�������Up�&��^Ӧ�����j8����۞�O��� ���d	t� ��C=T79$H���~^�ޱ.`������]����I�����4k�L-��F�<�}��p���(pHC�u40�g,M&���E�� �6���
q���{��JJ3�����V+�CH��u�Z;l @z.3Ne�-C=���?����J[�zeQ��A
׉�<T���J�R�Y�
������^;�-y�TVFb�|�K���Eb��ğ��y�e�$Ș�7��'��0���,��Aa���<���2��'��I��ah�/G6#�� э}G�o[6���&�D�ڄ����A9_lXvz�~LJ�0�P$Z��e߶\xY8�Qt�>њ����[z�;����B�,�8R����]N�A]��%��hT*�E��p���ŽY�͐���X�%����]"���b�Vw�ƺ�����u�LԦ,=:y��(MJSz{mv��'Җ����K�3�2ND<dr��Q��,��3��>��%v�~�R�PPE5���Q쾛F�=�*��B=Ro!0D���g1E��kM��ݯAt\$���.��ПY���P�����xJ<�w��.<�z]�Z���3X��\oƮ���_>��[{�
;=���:�|i���E�T/��_f��� ��e���-�)m�jO=�BY>\�0��i�=e���N�����%����0[��< � ��a���B��+k��	�C;+u��ϧ��0�@R���W槡����>t��:��vE\`k���(8a��6\,-M[�I�6�qCQ��ְz���9¢�a����n���5r��7���{"- ?Ɉ��A���}Q�4p�X&U�|�N�Ԟ��Gή:N��.վ8t���?�o�x���L}/d)���/��>� ��X��lo��j�߶Q�td�}iآ� {�ۆ(ZY*�DKU;�Gc5#������R�����^���`���Ier�LGz�C~��:�a��Ti!s�av�4��`���'��H�R݇�W)1N�p�2��V�\��3��5�*zl�I�s��pا�h&e5p�ƞ�7����G�Tz�E���j~ib�+V`��Q�ݤO�����e��/1*6N���=�j� ��r1�?Z�[>��D~��z	0͎�-�I>EO�+W$]��3;ߊ�����x�R�2�O�]��^�(+QcA�g�V���x(z�@<M�}����n��`��[����[i�;��-��I�Sn�; I2"'Ρ<���]��m����Q��th�^U�<�07�A�x��;X���MT����y��oإ���9��O��e�fl��i����O��(
8��rUz�\�L�<ٟ����֚_\��'#K��*W��g����UP��7I�?��P���5\�]���U��.RCh�5Ŀ2���2y;Zg�?a�D�1�8)v�H!o�J��Ok�y@⠠ePʊ��Z�n�tM���w�Uv�a�Gb p����,��"�:t0���l�_��gQNd���K~��$̗�Z.�ƍFB�/Xί8-���ݞ0��5�`��G�3}"�o��~� �~Ε]��c�\�MZ�O�Vf�}�(�-ȻX���H�Cfq�ya4P*g������*�ҋ��K���Ud���JZ&�p6�� �Ãr�V�R�聻s��쬍H�G���:0����n���a���k��\�T�{E��@�m�ԞaèV���d�b���F�k�]�W��.���|�OlD^��kF�[�==���$fՙUTd.�^�gt'D���n�h��7ǉ@F�sCq��*+hCBtb�,�(���� ƐD�ϻ��W�Z'��ag0�,c�I˝��F�!��H�5�%�u����X�ߞ�ï��l[6��Q�?���0�����u����h�d�j�e��-���K^��Q�>|t����/7&�u�!ƾ�t�ܕ����E+8�mJ��)� ೡN�
v7-��Jc�ͥ����eZ��V,����4���g��@dѴ��/��Ǐ�ۮc C��/�Z����h�^���@��ٓ��_��h�ؿi��tO�eHi��,�:��7���������P؊��ё�r�:&v���	? z��-��Կ��n��o\B�=�S]���!������4�G�INVeX�Hj�ƴ{߄ެ��V��z��Lx���᧳)#��^���Ge�]���6�|�:k'�"|RXﬥ�
*�0#����j@d�|�ɘ��,���0�i�Wí�5SƮR��{M�GѢY����IՄ��,�v�_�	�E$.G����ew- =1�@!b!W0W�����W�alr�B�=��T>5�i��a��O9�0L;��a��P� ;}>ġ�|,�:�F2�?���ğ)��-7��t ��0_�o�1z�������P �|���Z'�j�Ĩ��Mr� E5Y��+a� '_NX������\�d�!��U6�D׽0�8D�!�G��J=��t.!�|�;z��y�Od@}��D��A��-�+22�@�"�t�.�z"�Û��\���#n�;��,�d(Qa:b���\  �ƕ5��q��'r�eQ9c��a 1h�p�ۿ���� �ʦ�%���@���)�I?�h���"G�/N���
���V�P t%���E|4M9�{�J���0�#Q� ����Hr�%��wg���M�VS����|�k�l�o+��X>��U,��/�'�U:��� �k�T�k��أ�Wm�G�?�D��j�t�5��;�ѣ�52�9`�ͫ4�t��|�) ������w���l\Ҵm�U2�.\�M�����Y���o�O(����� ��?��v���*��}��\+L�S��N����Fj�(��8g�l;iE]�D�ap�
m�>�`<�#�m^i�� =@l�����w=����V���H�T�^�*�P�����OZ�I�q۹W���t��:#V��`C�~ �L,���,�F�D��p�M�2��߀Q����Pа쬌�;w�TJҘ�m7��\���d?r �(X�7�!��\E�?:ss���Y�*��(��9���G����o����������"[嫰�2�g@��Qp4�)�����[#S�ES�1�h]�Gr�"ۛY<H=RX���F����u�T-+��FN�Y�����"�]�S��L�H���("|]4J�� $��� �ds\H˞�j��S��9����T��:�mm��I ~���� ��N܂�sHd���=�kb��ϗP�dy����i
���, �,>ڢ,x�OX��n����5�5ePX��qȘ��Yb��{���e���
�r�����y�α�6���7�?vd�^�(.\�??�]��p�ۚ�y���]�b�ӂ����<�����d��h��N��L�,[Et}t_�g���P7A2�}�}(�1j�����_��n��o�Jg<���DX��}����|�$VX \+�Q��r����(l����]0a��Y�GJ���o�'�A|P��U3Ҙ��������ш�|�pH���Z��A��#��viUD��z��k�]a�^)ݣ����t�ꮠ�
��bj�I��o����+,���D�u�_Zhp@b�f���+4�ڇôR����XQ����s%�h�2��c�ﻠ�]ߊ���=^P���=���J�Lo%`�85}!���t������Na�������a|p����<�n����u��<mCYvo3���wE5	H��%��	�����Vw6�=�H�1s�ЉV��Gέ���R�_��)Uм�nz�^�(�e�p�6@y-���qud�K��8�P4��w�,Q�Mʶ��q��tB���Y�Ѫ��ڨ�k�� L��B]q��&�KT��W*� J�C�bS��`��G�s�hݣL-LA���?�Х�bSM�%���� 6-�U�uHz}��9Ҥ��Y�C�e[@��=�.�ZM��Z
P�Ⱦ`z�A����q��L�v��sM�����?m�q�?j�-v��;����<"��[�t��3����"���S�~���C�����8G���ƴ7]?D�з�B��3I�D��`�1F����V��� Y���r �O%��o���I�k��l"�f�&�lH���K%����Zq4��l��J����-	�Q}�Q�(���
��2��VI��c�J料s;�m8>a�_���F�#�"c�е9�m63���B�piN�ࠣ9|���~u}��	�y�IU�j���c�Ǹ�ct�G�M*7����h����*��������_L��8�^���3�������_�y*�Sˉ�Pz�����矧<��'8I^����!���ԝȈ:�%�Xk,��)5
A+q�\օ�r��FS)q``^�,8B�mA��3����=���lԡ�+�{" �>8u�It�<j|#v�'߶z�]�9�:�&.�7+��䜷��a��$���m��"G�
\Dx��A9�d���l�I��h`��o�`J�i1��8`��_y�XV�U��d4���X��Y���O�+0;�A�X����>�)Ȯ�M��͚�<x^�^�_�E�S��K�htA⻐gm0EX�E�����/bxe��!�l�$�1&L��Ӑl�B�@R�:Ö������R|S���7Y�!J=�D�WI��y�Lc_�_r�[�M�ꂕ.b��zY�?�k^ĭ���2ozGJo\r�-���_���4>�ѕG�G}�7i�C������q� fn��oO�.%�*�ÙNF���G�ؑ4��gOm�2J�X�Y>����P�R"OpƘ&�d�j������W���e���zq�K>0SP�x[�+\A\�y*�a	?A�����lp�z��� 2��{��0&��'sѪ��2%�d��?�,L5y-?M�m���'��P�����)�Z�C�Z���]��6.`10�Їʔ�C�J�\�f���R��+i�/B�鼰�8��5*u��$|��V��!`?QB]]�����[�K��%Y:?�5A=݆)v��~9H�݋�Y��	��C�qJ�/kCS�������C��vđf;�)p-�Ӧ�h���ݣw��κ*���F��̽q�Vq�� ��/��������O�B�Vr��|)�_0Ҽfy	mm(7Xz����LWݍ���F_�r����p)}�Q ���K���E_���R��9l�S2n5��(�����~�ƕ�H��^f��7s��L�!�D�R�bo63�*�^��?�&�"`�V��N�Jݾ�rA3ɮ=e����Ӑ�jR]���x/��oE�uh�l�ײ��i���$�rL~1\�`<=h;�e�C'R� �y|n�R"�F�p*<7D;����z��:<(b��?��������D�<����s	����8�[�
�?������j��)�2���ڈͧK�DZORջZ�a�y��~s�B��r8��v;�x��@�
��l����ܨ�r@[���7�d��$�2���-) ǧ�f�_�)��vc
�oQ��]+@/�g#6����� G��<V�Vt[ag#;�p�`����l<�$�I���������e^/PM��� 2�+�>d�߷�:щ}�G,:H��.��U���|b�����I%��
�~���sU��(�%l��W�G�q���2�.�V�����Ljz0r��L�q�J��ϒx����k�՚�J4n��?hB�
�z>mP14��6� |7���+R�S<hAg�}�HG��t$�e��,����eQ��p	�FF�8�(S��+s�t}�!�E���֛�nwKܭ��S���,�'�* ���ޒ������t��xळK��a�_�@��GG��qS�5��#�
h�9�Iq.���C���R&�j��
X'%pI��5�$�>���b��2p�x�E̞�-ἴE�:#S�_���(���Z�����/eH�:�q:6Ь#���t��ژ\4�M���S6=�c8��J��*��L�܉�ԐhC/����	�bꚃTB�(���^�Z/놘_�;qF����I跂��H���2W\�:}J��Jk�[<�%y�f2#P}��M�RO�%��Tέmh��Jy�;d+��{SP6_ˆ�ۼ��qlu���'��ag�q~HSd"O�eA��%[�u���4K[F�@��)�Y�7Z���g�7TU>�n,� �����&�f;��g�K
-�F���f�2��,H|ƣ��|;�j�ާ �J��=�32B�c�v�բFc��  �O[�-���z��Xd�n22G/�ai��Y"�Nbr���{A֚�X=��䕏.&Vz�).�ih\��6kъ�z���Fd�����&{G����
Q�+},l������k3 �ۘ����J�k�����b�#���x� ���wv�7�f�B,�W�{=�(���c+dn�/d�s0mz<A3 ʁ�w2��V�>q$D����x��&d�|u�B<��a��{l�q���,����A.8yG ��F?\8�'���g,�"��ާj�/0뱰A�gx�{��"+�5t�k5_H����@,��U�f�����-s�,���Щ���fu��	0��n���Uҋ�!���N�7�{3_Y����ʓ�%��͘]�8,'������� z,{Sʲ[r��a�֌1
�p�_L����p'�x�K��2/��΅, �(\�&׳���"+`[�s����I2�Å���!ŀ��f�RgHu(T�i��b9'��֗��hm����q��{�����qO$.��\����((�ܟY;��Z�9ch��*sf�:�#n {��.F�m&�����Л�����"�Y��pv�i�'�j���b,�	�_�n�\f �q��A���!jo���J#�V�v�i
��/, r`�V�DXc�o�d�� ~���N�b��\�d�ty�f�pwc�����s��?�c��7�o6�'��x4�/0��%�:�� ʮ��E�.$�/�x��Em�2����}�謧�j@�\��폯�t���m%�I!�Wʩ�--�y�yx�@�XbA��D��L�J5*�C`�`3��f�����`P-4��_�	�T�:d��n��$ ��C�Z�&D<�(�j~#���ta��
��u���j���KOڵ!�x�y��	��M��M?apba&<���Y���-
Mh�*ەZq�?�v0h��'���޸rsKi�6�S
�.nh	E�~�C�&M}�ϭ^G��g��u1�xk�$��,_k(A�H浺��V����"d��b�8���T/��J�$���.x5�5 n�/W�W��aiKoc}�'5�+&���A.��l��Ǩ0R��޽Gtl�Rl{=���/�$�d���l��0�.��S��-��&	�3	�٩'$׻�b$n�������ٰ���Sƽ�����
�r}c�*�M��� ��Bc�[Y�-P��i�@�^DJnT1��OT�:�d�z�W���F�~i�br;�U�8���{;4d=�cа�w-}�m��(�2CE�W(�0�Kx����˓�F�&�����f.����;��\�k����D�O^�Ĭ��8�� U�Z뙻Z�_�6Z�d���������#�5�(cM�$`AI"���
D�uN5zR��6<i���'l'1� �֠5Nm���U���?W�$ycYS�lߴ�5�Y�W��#�Y�[bHZ��3��t0��6�c�W��<Mu"$��y�/m9�z�6������7ڎ�Ĵ��iQX����EZPCZq�&��ư�_�����P��l7K~��C2�86�#����}R�;[��R_bX��/uъ*"�F��y�Q�p4"��N�u��>���%���WQ|�����Wg(��s ')0�+�{&��΂Q^�����T�v��-d��Ő	��br]��z���n�|��~r��<t��pS���I�뙺Κ��.��F&�n����W��J�XLP�K�5�Q*�v�#����������W�H I�HQdA$�{f�ב�S�S�����ÂƬf  �V�\�> ʉׯ�eOV��	�爙�=K[��h�J�O�"����?�en��h��jhu���A࠰�\�!C*d�r���yo\M��#����/W��͡pl^�A%Ǝ�1a̡��vN�H�%����c[�x~��`�S3�g2%�^t�(�@ﴯ�]���T,�*Ho�����5ξ\���
103�g֧���@����m�n)�Թ���)6l�a�-L������\�GEL����sn�beO�]�ٔ���(�$�m�+H�b���MD��@4|�a�0��\3*m`2�[�QuT�sT��<�h���m|��Ң�Wl�Z�ܬ��2v��?Vg.aZhg�{�i���dJ�/�����/Ƣ��Pj��(��V�O񄖥�CɺW��lf�Hv�!]���;}�&�_V�6E�Ps_gB_Um��jP��i�g�g�
O�Wݿ}��xZ��pK[�X�"/�J��Y�q�Ҥ��a�ۋ�P:`�Muxؙ]�)����'J4-Mξ%J��t��P�H&�
���F��=I�0k�^z����Й;�����n���\K�գ�V�����]$*һ���g���n!g3O٪�l@� ��W��+��&�_"�1>�V)d�d7S"qO��	������GF "���nP����w?b��[P���\.(w��c5��d��Ѣ��g�eV̧j����ti�LV��/&��c:�����ГyX
���2CG�^ �8��p����U�D��)Nf#V��O��Hz����M����U�h-��L���'W7��گbU�%�v�p�l�j��j��u����Bf�އAH[" ���$���<��Qc�fxI��H~��;#�%���I$f�gP�C�5���wȰxm��kq!�uש��Z��嚞��f��e;��qֆ͝��Kz?jD��lZ���v:}3��P�h�Et�\��$���;J���|XF�& �lb�`��	�s7�==��O4���H�a[鲳H��:�j��,��,嫩<��  %�=Mdm�a�0�6�n� �4���߫�f��k�$�Y>�F\�~���t�t����V��7�2�78j�-�l#��|�W䙚�	�$\�d��n���7����]�k��{z�k�����5 ��_N �Y׆O�N��/��S��^27�YH���R��� uCo�R'\;��T!0�ES&Z>��a�0���|����٢y4�<	��ݬ�y��;���ԣ�佄���KB��)����\��=�h���8�k��R����B�@XW~��.G�W(f�wr�N�OէTY�n�ʻ�(�y�y�٦�{�ƃ��>3�qfu��̬9��?`��7w�臵!��]�9 !0������K���{��	Ӕ̉53�dl���5�LHsE���7��s����ݰ1���)���(#�>��5��q�-X�=%��2��U/ո���� d�x�׆�~-v����<cg���-�gL��ʵn����ơ5<�^�w�HF��\���
�������'F�~u�z���٧g���Wۻ6
��}#��_鷾������2XÁ4�Փ��g���ƣ7W�'��X4�Zb���9j����-�j�.��
Ē-��h�{R�W=��3�{G{�ճ�x�]��(<�}_�I�uOr�"�Or�_��3Ӏ|�H�/��#%$M�S�/T��*�qn;���iƘv���b��l�F�橨r쏷$��.�+.R��Q5Z&h�:�;�q�ã��Y�E����A�����	��&>��D��;H�rӑϮ3y.����'֒�긷��y�������@%�|���}e��H�TE���TQ�3$�����_ ��E��{�`N�
�yܩ^sK~��x��	��ci�4�̀�t���+\��ｐ���2�Ɖ�"GN.�G�mv��5>M_�(���t��c�T�i�HI^0�b�-�t��{���3[��3|Aanέ��*�!���?
$�@�H;��Z#�����t�m�O�ԯ���������L���6�c��tY�E�T_dL/�Dz>�.��Ú�0��;���tj��:���B,�*ʶ�����.�C%@%=���d)����Ce�D!��$�`c:��%;�h����h�~�����K��|���z@⸍+�<6��_%EE���ͻ��)R��d�!�Z�JN�ob����5��H�YX(�!����65�w��~)���'����P�e�۞"0��f^�ؖK)���Q��R�
aJ�+,K��rp#�''2���(5jc�rUq�V야�Sd桠8�G�M���.1�/w�2� ��k���
"D��4��F[�%��u�FM�I���*��F�I78��_�P}<7o\A���L��(H���=�?����X�z�y_�"#��9b�?��X6=f���ud�A��!������
�5��r���O�����������ۺӭ*��̼i4�~�-q�1u��� �:���Q��FY��g�a�m<�aB4*�W��B�D�r����;�z�2�>�rX������P��f�������e2��c�y�a�
Ny~ߗ2�w��<��j��&pk4��7Ca[���3C��Р���G�j,4V��ʀݓ��>�gYj���:q֥��0HyzMvc��]�@Uk���V�������~��6\�n0Z���L��|��ZIh��z�|1�cZ��+#Dpv��,�F���� �H.~2q�����8�{
r|�2l�]�?^�ހ��V��̚@G=�����;nv�#Ȉ�po3[bX��񓕦�Rv8�ݺ�d�����z{�������J;x����$�|_�dR�>dZ�J=���r�-<KPbf�� ux���}�З��Ķ���k�V0��ю�Gc�����hKB�'1;Mԛ���;{���>s�\��y�I�;&]���*pw�ߐ3��0�Q߭nb�;��K^���B��p�<�e͙����"@�Y�"g���Q��|(��©�j�%���ʻ�R�� Q��5+ꂳ�tɇK���q�̛N ��E9k��*�fj����idM����V���X��!o��3�|��8A�]�D�wb��t+��䪸�P���U�r�{�!�y6��!e�P�qo*�0hw��{���TZ�1rdi�Qӌ���o�-���Kc�/��@���" W���QAee� �Q��S�\�o�r�O�.�[��}$�`$���1{1硐�L��Vx�w� ��ԩU��?�Rs�s��� Y��>�.�]l�UWE֫P+��F�( Q��z�Aq���=�| n%M(f�@�.?k	]�"Z�HT���f��ir�S�s�;���6�LX����l���g6I��m-G��:r�6�r/��'�)���Y�C]�����sX���e��	t��_��|�T��J<��(6�Kma;� :h��ײ�f-2��*�!㌌�C�z)�',���m߼!�-�w���1{��a����D,�?
�e�S�\���c�jK�4̠������7�\N��������k�O�w���ՆĲ�q?Q��a��T� ��#,� ͉�EP�s��t�fb�*�9�m�!� �k�A�Z������Mu�/�҉�0�H~.!,u�K�����]�77�
�Ե!�Nl8G��1C�d�&F�߯1�t�'*��qu^�%���Q�!N[W�7�Z�1�V[���y!yB������	<c�Kl�̻�վ�CKaF�5�v���zB}Nr�_����/�E6ۢ~^�s�h,�u:Y�	ln�t1YU��!av<U/��&"_�'��G ����9�%<�X��G����b����L�!K��Gm�$y�"�iK���PO��X���:�G����U��h6��Ւ�� �D6�S
��j4rYo��C3��K�ll`�8Z[�+�m�1��ѧ`���>�n����|����.�+0�:�v�b3���L�Ϭ?3]>���珛���%����˽�;H?J�[B�E���q\�����Q�>�pۤ��'s7���cc�.)�ŕ�O���������x�%Xa��S͝�7��`&'��8���Y6{�r�5�t��R�?h���o��ʃ�����B��2x��)k���`#{�o h����A��7�M.����T#�P�\��,l0Fg��ސ�����:�WJ�� #U�!$�� �Ϋ�­E��V�T�@��p��T �I�3i�G�=-��Ck�͊�rG:�h�.*�{�&z��R�..t��o��` �ǂ(���/i�`� �+�6.Jg��LE)SY��p��v]��җm�� ��<�(j���}[�>��ύ�TI�I����Y�_M��7�2�$�t�N�c"�veB�$��GQ'��h�Y.��eM:I
h�aę?��ҸaMo��Nn���t=Ejs�2�܍߷���e��|��b�YD̂�I[�i�T�od�o�A�c�_2�ă|�n�����JoS���Μ�v��ɝ�c��Z�KC�g-����/L��.�&̑�6���ƪ�*����r�@r��Q}��;�<\���xΕV����ZR

Q�| b+��(:dv�K�(jʇ������}�����}�{m�տ��O!__3U��3t
y)�nD��̥����Z��Sfs����۳M��Z�-��½G��5�Me�a��Y�?W�~QB"�s��/� [�Pk����ʂV��Sw��`��{�M|ß?ic}��˵�z�kke�5�Uj\_xM~�9�+�Ԛ���j�=S:���f���`��_���]��[@>|@�h*�����)0�2��������|���K檕�!�lÖl�M���;d+1 @|i��*�D����2�o�P�ˬ�"��;{���8�s�.b��h���ub��Z���}[w�8���ˏVi����V8���5���L�-߫� <g^��5����*�!�7�	�l�YEA#$�[�� ������������Ř���?O�e-������Q$3]��Ii+l}E;��҂|���t�b���Ū�E����X���dHE�Z�����M50,�e�|��-Ռ�%��1��˪'^?��fd��\�G��31bt�>�9ǀ�/Atc�[�/SK�ˆ3�����vA���?�A�İ��~Q3Dz��mL�������w*NH0v}���6�2��(��E ;<�Y��Su���ˈ��Z�ۨ�Auu
�	-c"Wٷ�C�1�V1�4"��bE�$����Қ��K�*Z��*�na*#˙O�ڋ)O�\�U�x#&K�;8RF��hZ��ņ�g[w�H���򼰅;U�v�A��w��MA�fF��SX��e�G��6:.�6��<���lz �s_�������j����լq�=�<t���l�3�ԯᓫ�@�l�Z��ٙə5�{nӔ�R����������7Q��?
�yj�~��[!�BZ��{�MH>ߗ����U�S�4,
���T
����'�!4��cq!� ]��_9���X�ǿ�,J�3�V���[���N����/èDt�g�\�>9��$	c��=���:��;[��u�]�C��j�)�����b06o����	`m/�=���� �,�\�y?�0�1�鑚eRX(�Vk6��/�����8b
�H��z���+edP#k�m���Z�ȥ߹��tW,����01|��� �Sdc��4����E�\���Nʤ�S�/���bb�����~1ɮ�v:-<K?X]T���/m�ݍM�\�|�m �̥�/g�0&���s�D��e�9���y�u�^�Yml�ߓ/�����G*��N�66r�d.^�tF����=ìHʭ�q�l	jH Ï@�1�Iu�"���7M���9s7�����V�e�&�9�?��]�-����\9%{��Ҡ��J�7��@�JAEQ��CH?�طRu��O��xܖ^��Z�:�zq�o?�O��}��MQe��p�}=����kZ�-�?�V���ě�eCd�'�i0'a8vB������/�)��#�������=�&�>1^^E{V�mA���������q�[���Y�jA[���(F�E�Ad`*��E�$A��2�����z�pr���|��O�	�� �r����CHgL���4�؇,I�7n���C�o�y���o�C
A������1�@�M��ٶ�t�wG�R���[_���@oaTZ@�s��j�i����[��ԩm�l՘�ɋb��L��6Ўsk�������.�i_g�_����׷�kT�x:G�ݶ�z��,9AGʍ]�9ю��:<���բ����l�qd��o��%wuts^�v�J�>���q�b	Ⱥ�ib}?���S���$� ��r/Zl.��)A;PW������o� �H��$hsنeD8����~�B�^��ߖ�̰:�ԗ�̰���h~iL}*ޛH�5�D���4���x�UR��V��>�m.�S�3Se����^����9)�:]�����~n���_��@j���� �����TK�l��t�HN14M�VF'QI�"y�%kul`w���8����܇	������{�)���H�}��C�W�,�ї@V���oiC�c��p7���G�KV$�GXP��P�$+2c.��S��ҏ��2,��� I {���ԛ,���d,�맩'�8OE0�C��2>K�օ�W�U���������K&̈lN�8e�
j��}&�#@1��?Z���J��C$����5ـ���X��|�ba//�!곾.��ia]��k.�+P�oPf;.�[Uk|+6�!��[��ߛ�2�?�GZW�j����3o���lm�ƭ�djk5�ԡ�[��?�ظD{;^ȭ�ptKd�n%�lIv������`����$�x��qn�^���fdG�۔�rEi�Wg|�%n������
�#�~�Λ9h�:�ͫ��e۱K��i)�"��mLZ���ܢ팋>�U1ƅ�XNj?[qq=�z�Gɸ9g�5N��Ā3���%J�bV�	����a�T����e��.B��12lЛ8=��$[(ߟc$�[�=����8�.�Ag�������\O��b��Rۑ�9��*�"v�� �d��~��)L�$�t$�~�"���hT>V�7��Y#(%AP�L�t��7GȎ�C�3|�f��`3[��_i��>8�0�8@�5r�:&�Cy)��b՛�\ȃM���V���b���Kϭ`�I��N0�����iVC�kQ$���0�Y�l����.e)D[�f����2>��S��4G��{:��l�'F��Y���I�����£�J��a��b�|�v��9U�ˠ��gRA�qBQ��6�4�$`��0U9�"$����^nT�IO��\6�X�@�E��W��>�=Y}3޷��/��3��1UHC�ᶦs1ܯ"���������趨$��횥[!�ʬ�'��GE����l�%$�?�R1�
�@���0�����#Sx�vv�i�����~ȗ��Ԧ��$�0��%˹�E��J?��12m/0�q�~��?,E���f�)�@��dWoZ�����/{�W1)�
n�õ�2�+�,�!m:U��Z�#��ʑ_���.@6�C[J?��ڞެN�n(��a�ee�*�I��
xT�3����Z��Яf�K,Ҏ����nFHj�����6�g���e����S.�+IEM*L�?�i����֠¼�赮b���	rhofarC_#K$5���A�M_����o��I�$(�v���[�9 "�+w�ي�n>�z�C���ƨ�L��mfP�!+���?�T�(�W�����4A:��Z	[��^��#�[rV�<@x���$6�z��l�M��p
qR�3Q��	�j��C�~�pY���y�Z��v���kC��N�a]�ߵ���`��"��X]V���w�m���'�v���)uZT��@��ۏ%��t���@9����
�k?���N�TWQ�����,���b���|fLp�Yӥ�&~"�S.�?���%��C�;Y�+���Q��&?Y��e��Hq�n�O>���N�J����H�r���������1ѩ8�!%��,���*����%�=��Mm��{q\�AgW�1�*������Li��o*�d�Y&�e��7���d�ܞ�_�q�x�jzy"�~�m?{gZmK� 㾅�Ԕ"���b��}u.?�9?����|=z<M��C����{�<�S�t ����ת���^�]������M[��'ɫUܼ�Dd�Qy�#�_��f�]������w���m��+4Nx'�_;���7� i��0z�.9��.���՟T̩r����˝�h�8ax�8�� �	8� ��2�n�������,Lf%�hf��K��1U���j��lV�ƣVz��D��P�����i�W/�ߑ��'��_T��<�3�{֓]�iO��]���C��1Uq�|���!��;�8\B�*������5�c�N.^�|�'B�꜀vM���ڕ��btOk��?my%�ߔ�7%�����%���"����`?�	2"(e/Nn��1&�/�wΙn>Ay:�uīQ�}9R�љ�g1�+`��S�C><O������CG���fk�4|��SF~84��z)m�i)�z���w@���0��?�Nz��� ����yln�p8Ms#�6�6�xr��(���b���X�h���Ш��}�5�~���@St���̟Z�
g&�h$ o}?M��0�D(i�`+�vK�m��65��6�=4�"�k�U\�����~b?���+�@>�H���:��:�����T�:�`.��A����Ygv�^.I�=@�7:�H���p4ᅌ��-R�l�A>L~Y�}x��PśX��/��eJ� ������p��,����G�/��ZRxD�8�z�nYO8qCFX���Ye��C���W�<\��79EV	�ԇ�5 
�˴-,��[�
�*j��|r����oR�|,ٗxn����Q	:�W�*��?gd)�~T�Dq��M���g�t�p��#F㳫���ڤ�� �1M�����Q	y��:Ԗ��)����\�H.�x�j?G��Z��{�"�}���)�E��E�P5�>Џ�O���Nt�;~�t��C�h�S��úb߳���B}Lu�XK�`��u�O��P����#A�����:G�^k�o{&��\���we�M��ȿF����1)�
���gO�#Q�t�ӂ��������I���Hp��u���-��YjL�ΊGT�H�C���K���'�%��@-��*��7����t(}�ח��DY����ff�����FM����N3ő�SP�_�Ep�\w�z��ye�j�C�@��H%R.A��ji���=KVf��oYu6uBк ��RMy'
��m5s��#�3v5�Z+���IPr#U��]�# �H�]B3�ߝwn7�^�q�(��]'�|��E�s=���X��v�/�7So��!O���O�o�'߃!��{���N�I�����"��E�%��Q�
����&�ޜ���,tY��탰����Dܦ����:.�+l��m�T��Q&�A������9Nƺh��㰋k]���bv�>����8�If��u�?�����J�e�q�T��)xm:�t� 1��^Apщ����1-1���aDRM+��*�aF̼H��f���/�8�$J�������n�F5���Z
�,��ND8�����"��c�"���3� �D:e�j��hy9��(v�\��PAx�����|��~��oy����N��rQ�M�$�VWz����+�^��f"K`�#�snΝX�A$#�C| [�"����-�+zU%�����m��̟y�B^�X'�yo���Ë�qM=����?�.�����C���b��3���E?��o�쬶��:�̢�O�;�HR*E����ؠ8�P���ek+�k�íN�Y2��9������g�'�T�-��7�	���(h��.6BKW�&�мkIjKl���ŗ�g�A+_���,��N
d`�{�+*��w;�������<�E�����(���F��`��H]+��$�ܖ����`�~�3I�D��(+��y���2x��_����	�.
7����$�0���N���Q+&�,D��sܡ�E�g�C�Gwtzl����6�0��T�c��j,���|z֜�
T�&�Y�I��vY�9(mx�#n�a;� *p��3��Ҟb�ҏ"�ARFY�g�B�^�������4�����ͯqH�)V6a��[���T}cK�1$L�y�k^��A͟��~�cܫicx�]��*Km?�O�	���Cb�&�LC�~�b���1㱒r��d"��=��ۛʘ���i���$��T�"�PD勓4�m�irh�Rx��Ŗ'L�M����>}ʍ
��hTǫ�q9������\I���I6�Qz= ���jݥ�&֡?'q��,O�ߎ8�\�jR"���1Њ�O�>����O�9�j�l{��ҫ=lXc�{�z�x����%&���A�t�T+�C(mW��P6\�X�s �'��HF=p��%��w�I4�n��l2I��1���]�썚n�
�*���]A�1Ӿ�kŖ�Cz"�z�x�Nwb>��xg=j���,����~,;qO@���2YH�|�!��d`u�l���Soò{���������M%� <��z��-m��[5� �ZF{p��B�ڕz	'�	]�ǘ(��Y6��:н�8�Lg�9����+޾�և��Hɘ_NW���� �',bd�
��a���^$Wo��Ve��Qhʓ�;:�I���y�#��(i�)O�[{�?݈S��wУ
�B����@zk����t�|U���y��m��@4c���6(���(�X�m��2p�
�������y)�-+�%��
/d��������)�ps7d/�I|`U��ȫ����hS�V�*d�E�Ia�k�sW���sU� �#���;�_)$3��uuHђ����nq���V��6
c���3����1ǸtpU�O��pv�RIJÇ`z�V�(���g&C�z/������J#��Ֆ��de��.���ؤ���*;x�|�R�$�;5�h�Z-)I�;�Â� J�t(&2&ȗS�A5k�+�tqC6�Tf�]�#	��2��"kX�"{&}��g��.p�W18�(�Z���eU�7Г���,`�E�!*�C@��c�[I��_���Fg�̈́Ǆ��hS��!��1�?�D�XY�����T�gظ�Q���)X� .�:�,�.�6��o9w^��Z�5�d(E�7��&�D�v��#O4�rh-H����\�a������$�ڲv�4�1�V���1�
��f��j@�k�y�?�X�s�4��\oo��~�خ48�r^pD�(��
&��3`��NC,г�
L����$h:����0D)#�A
�RcP7:�q��?���%��B�-�a 	hQ�����D6�Ѳ�H�玜������{c��V9c/�Ť �:��q>/���bˁ!J��J�;�n�ܚ���X���o_��_���T�;�bs'�Ƭ�I�z������F�O�&A�� |j��7��S���Oh��5ڢB��X߮n�Ź9p��- O鰺w�˸��v���w�S��#����^��01NC-�ɕ|)\����z
O8C@�#��Pƕ��v�'��\�K�0���X�f���4]�'�nWl�h;�z�$y��E}��Ä����)-��+e������d|��Uz*�JR�d3��7���x�����F�Uj�카cŽv�p=��Ɉ��M�\�c���h�yC��9�=��;���q)�!�7A�@sLfhv�5��Oo�;��֌�8OS���$��3o��xK�ޙ`�&FK��&�~�t�+C��oX.��j`����	��wo���,Xx L�f�8��\��Zfܽ����s����7�v��F!�n�_sv5�&�%'�Q�h�VXÐ�����v��������}���!���/��?'T�-_y�p�p�_�$wie}���}M�(B�x� еP�R1g*��ρz��6�ZV�Ag��H0Q��Q!��T�;8f|8�)����q(���S����_K0"ȥ�2Z�3�U��+��|�y6��������{<��H��i�\�'.P�P� ��(牎'��ㅞ���Y�\ت��ӿ�"r	O����Jϡ�'.�yA"`tm��g{�����L���\!�O�����k��MNۂ�M�nOGo2�V��7�2�V#Q�?.s 4�f���x��$��[�bmp�#��+���>f(L��ڹ"~�,q����~�Y I������VN�Ɣ�k��ZΒ�8��D�����@���S��}Ҷ�[ў��¨���"4��&`J3��W��8�H��;q��0��I6�[?�L[$�.�7+�9)چ��73&$��b�_3`��[�G��#4�׬u"^������.�m)�q]�{�<���߫A�񌅔�3�ʄ]���S-��?)Y�4�uo�NAM^7�ktPJ�4l���7J�$��5��)��y�v";������]v�׽�0��r�
��x_�b��9)���!��yD�އc�^�}�p�R3f��ޠF��n��F&��Γ��4nl:�C�4��}�l���Ԏ��=F��8����X!��QډvWp�nZ�����_~����JpƮ$�0����i
G5Nm�����̠Q�'eM��K���O�\y�GS���*�⊑o'k��(�`eQg�c�O����v���~CD��n��.s�_��Pa�ΩH5g=�4�M�G��5�E�D��Eц�Z�m�d��	�]C�b��Ѻ<���<^\V{�����4L�ŗ0����b�T��������8�B*࣪�M���GXY��B�*��0�:iP���o���>7���wu�U�I���`�ᘸ�7�����47�p�zH���,'7U��š��A?i�e8��Y]`X������+�V�c'�⩪�xGO���>���]lH`䷯�TCH	�"˲��8��.E�!��t&��5�V:���L������s��N�@-/pD��3-�Z��+}t"e��L�U��1[܍�@���)n�M�HIt���dI��P!(?9��u8�	\�mar{��	�3��=}E�GV��� ��sS�XүC8l,ДA��&▱Mkkl4��E���}�H��@"ۡQR�DP�>5�@��^1�p�26�����\�T�C�_y��#[��?^�ʅUU�zQ蟀�h%�A�9��	]�*�dyJ�y64iE�|��\�;���rhe$P�h)�_��������?�;0�O~u��>�LT��>I`�
%8`Uc���A?9�?Y�3��X>b��Wja�E�ߪ�Ʋ2�a��# 7G���x�*� ���6#������d�<*�u*�����٦4l�ۯ�[���ޔyIv�� z���n!�� g	�[5�!�,}���΄�����o����
�ߖ�c~!V-֧�3�k���*�kQ�ٻ�UNJ����x>��S�0�p�4Q�m��i0Z�C����Ds��Y
h������Z�;��>�65#�kݲЋ�����R!W6�hɓ;�����y91��G���5�2���l�30��BL���Q�8�7y�m��l�Zـ~��u�/��=%�"�$��^V��?	 ��ˉ���:�ևP%�D&�JE��TK=VOQ��N����o���AV�/���œgGy��oo6g{�7idG��������e"�T�o�x:w@�,v*�m��D���f�n�hn~l^�3.�f�&�(`O?d��5�����>�$��������J�D�l�ħ��$9�0�2p������{�
1�Vvm��#Q�YLAF+�%����0zN�ߏ��Y�е��! tN h Ԇ`v���0�x|�$�{Gn2ر�MK0�
]��ĵd��*��j���^�z׷.M�&2�+1׍e���`��u<P�o����lt=��ږ�ϫ�_���$G\�m���F��6pN�߈v���4�#_�N�n�в�b?$	U���4p��a��"#rZ�hq9z
n���ȤM$_�-�ʒH&��(1F k�����j��j$� mrx79�MB���&̿���H��r���Ȑi��P9z{�R�l
kp_3�O� (EbȤܐnpR4�T��ĐvM��^�G�
��+v���>����F�����06K��%���q���h9"��(we�qsx��"�\w��{�=�l���j�EQ��F�8(�����]�_���k��=�����K֦���_��(�l*qVI?n�����F�db�l���,��<��N�����m����y�l�~�<�e`�{wlz�A�9�F�:��W���LMKi��S�k�( --��Ϋ��jZ�3kf�w죆��ř��=��`& ��/�����d��25C+����z!]�2� x�q���ʞ�;����)��ݢ�q��`����j�#��,i�]�t9φ�~=�,��BN�U�!���叶/5�h�Y�v�!����(4½H"j�V��n+ʩ�r��S�xQ+v@ю���5�?Y����_�M@����4�\d�mT�.d����:������(Z��4�nDv/ͩ�c��L�\K�G��b�)��+|��������E�t����#�~�k�
��􎦸t��H��*:%�y��@?�sĕ]�x��,f�I�e �j��C���e�Դ+r�G�͸2��ա<�p!=`j?�R����~�X�ЛML@J%�T �x̬s^<KR��upR>=R>{�c����ל��g���bV찍��e��ʖg)3ȶ�p#�7ُ�h�t����+�������ސl���20/�~�Z)�)��2���n�qױ�ei�)��?�ާ���n��_]�
��3�����T&�꽑� �.>H�y��$/�Fl�����F����/"uTH���ӌ�F�r�e�7�E$9�$�H���Â8�\����<VDgQ f�p{]���+��wл�6!���o��$�L�GXϥaĶ�X�j`��M�̻u��<���`B�ؙ��˵Ju�X #L�5;���d:�aj)�U�Q@lk����k��&��lk�L�C,��qQ2c�s�� �B�b�U� Z&ә��X��e��+\�@K�Χ�k(�!�ڹƯ��\|����� q7FJM�f ��ҿ��n��Ȝ.�K�rH1�k��c���1*W�SUjo�gRO���U��~[���~#��gF����%쥿r%ǿ�7�d6b[#�*O� o;b����l�I�|DIR��GM�8
�M%����/�B��5m�RÏ6q����Lc��p��O|�gm�����F�&�0QA��
�U7j�F�iD�������]�Y��B��)��ӀRT�M�OG Bד�t/f>�'3a���b�+�oү��-kG ��uLQ�m�B�����-��X�6��\����I�C�J"�i7 ��$:�d�{��tg�R�g=;=E���?�!6yF���b�7Ȩ�z	a,,C��rv�@q����'���@
=��شYM�C���G��!(�E�vY���r��(iUʜ��?-��v�s��� O5g:��W�i<��{TA#H��#�<���G��*uP(F?�x�x�ӊ3ٙ�`I�����7�fm�0z�5����9uB���?�PDXLoͲ��:ܗ�9=8z�፤��42v@ց��0��0�Ө�:NZ9mc/��6�^}>5���CHj�R�:+c^���_�s�s~�?�3�ګ�p�od��)����������=�s�Pn��`H���F��~�#�C�pQHM�E9�.�ŅGWCozޏ��=㒄�Z�1�Ѥ��|�c;��u[%x\�-�r釋����=Q�;����=p�u�t��܃,�������5OlV�kG%����f	��m�3Ƹ�^�ٻ��ѳ��lCSbnTԬ�������_,��[��$<dg�:���S֫�.�ܾ(y�t��r�qĦ=�|���2����o�u��0��6˜E�.���}u��}���e���|���G�c�h{���f7�Rxq8�p���ucy|2���6�#3)ĥ� �N,���2����ZlÑG~���e{z�;�b�՘�x�;������!�EI+�N��� ��f��+��Z����*���x�=!�KA�A�y�� x��0�����S>�7��c��K�m���O�2�%#�@ϓY����\4I,4��XB@��#�����r��%u-F�}��.Nz��9b8B���d<�
�"�(�a[Y&)/���"�������@瀴l��UBV����N�Q_�b4G <7�)��4����
�x<X�<[�Fa<�3��*ayl�5�5N��Zv����N� H�������"�77d(@q�<B#4��o�q0�j �[y� ����6x2+�s�~&�Cz88�tm�'>D:���c7@~���ܢT�Y��܊�}AX���\R�����I7p�A��������!pm�ْ㫮 ���9��s�p̾�@Nj�^�$":�I9x�D�h��,���J��!m�t�X�xF������h�F������7��?o����}�GW�^{O�������f�0� O,:{y��w�
�\��O�GO��h�,�|��h	$9p.͟�0LQ.W��P��)�(�� �Ν"�����<M��ܹt��CT�]�<�]�\�^������|킂;	�?H\XtF�Lh�q
�sN� �ii|�fқY�W�T��$�:��f���j�`����׏�lŨj���|o��Z�|�&��r�p�
�r��M��귇�@���&FH%"�y�%��ʗ`���^]�&�������5u�/��{j��O�Ր{4�'��A1(��t�Mbj��Ims�ߵ,��o�2`{`�?�6Ȫ��O}cŰ"��D�b^�� @t�fW6"�{�$��׆r���ji��|\>~bR��J�^���^oS����2G�V���\$(�:�zѻ�׈� �F�͂�cvU����ʺr� ���a�P<08�m��<�
dh]�'�*y��ƺA���.��1�=I���*lN	&Z����~�Vh��@ALy���Fȓ��tќUV��q!!t4/b��u`K�C�]���j��'��-��L'7��������Y)=$����������$��P� UA�p�&�������g�ȵ�M:�?�X��%"���� S�s떭fA#��k���M��^�%�aG.Z$-�����'��&7Tf/?,A�10��U�FqCz/�4b3�`|g������40�oxx�Y�A�s��X��(�'���9��N�h�l�>	����l1h����9���_�p
�Hגv�9�GԔ�7��I�	�����cj?�{in!��a<3��;�z���<Y>��ti7��OX8nL$�)�t�Z1	�c��{�Wp-�]�T��v�{ætv�_�\?k��������v!�*�Z2p����T���������Y�th��;��@J$��)cg5{O�Z�Z�O�C�
c����^���1%I���h=�h-� �H�[���(F����gY��R��y�z�a�z��&�;���g��l�& �1�u���u��Q�0�s5�����oͅ��g?yg�G���ϏbZ�b��*�����M3�R�1�%ǀ����W��$�.ΥW54�*��p'�F2�.�jN�C;��X�\�Z{�h\��LF&bQ�1�zb��k�k�����i�k�U��w;���V#�$x�bN[.*��*�u&�m�|�=��)}oٽҜW ���?�[�$����XV��H��qQ�4�0k^vG�W��(gI�Afa;���Μ���cT���o�*���F�U�1ML>J,�C��:�b���Vʆ��@2k�ct��a�޵�wZ�P��1�����0	r��]?o�t>3|C����&iXm�->5j(J�3'��*5jh~tn&�
I�@�/�xD����9Ŀ7��.9U���/�Pj���3@�T]�Bs���[7�B;����o!�<�X�Q�	�7�Y�Oc�:\��HO\o�ے ����o������C� �`,̿��]#U������%9}n��>^L톮O��
���-5\~��W%$�,�@�}�������6%&����a�-�YO�J���L��������B�o�(��T��W[H����Ұj68��8]ئ[d�\�)`PU�a���E�訙J����6�Gm�-r#�������x��h��^�:T�FhW���e�021	��w6w��@_K�?��KQФ9�P#S�I�􋦩"$���A�)-���%՞/����S�T����'rAJ.�6�b���qF�Ɖ]$?��'���(
��g�sc�����Fn+mBK\`K(\����oVQ�oQ�%�o[�!�]����	���$��	�Q.��h=GQ�,�|�Wd��d4rfjѵ��F���4�S��o������Y��
7h*�b�l h2Ǡ/,�3��p�&�#��+���6�+�^jS��h�%<w���C�iy���uP"}L���g]O�]Ч���e-<(�%��#P� P���
�s.v�Y^jo�������T?��=3�&�~̽��ɶ��l�G��[Aʣ��eu\��*�"�kIB��y�����?cX�B(�צ�o\���t iR]y�n5%��jf��\D\�{�?Y3M�A�>��:��3��/?�h2�&���]���b3�OY���b�ŝ%d���?�ԩ/��r)tP�lS�ۉ�Wvz���muN���z��$L�H͚iWEǃ��h	���CE|.Km�m�Z�U@K�/��'��{�ε@1�>�+f�pI�?	��}{B=��3��2oSͼI'Ǧ����Cc/D�:Qo2�i��]���O�솮6��%_؉��dL~�+@��C����8g�DLD�=ۛ8:���������So�+�`�+���y�#���1����/�3�1 ����q��`��:jV�+QLK�Z$�Z6M�K��L��Է,�ΰ�c&z0��)ґ��9n���P�ŧjVH�u��Ȟ�<Q$s���h��)8��;����c���[�*����8�'*�v��<#�8�ɻ�X��� ��r�/��{s7��W�� g|����Ⱥh8��@1�k��̔/�w�m(<N�#����w�R6;<���e�{��ݕ�<���mS�Yֹ.���@����|4��΄��.t�(�����|���C��������� ��8׀!�v�:�>�i�ҫ��D�P�����s
8X�mw*��e�2�0�1�g}�D�[[B^$�}��A��'�'�\`ZA׾��H\��H�[ٽ6�i"%��f�R	^-�gj�T..'�dX%_�N��+/Q7����[��˯I�56���7D��^�H辪�TU]��$���%��)�i>�3h���+i��7K���*F�nű��2;R� ��^NX��p��D����&<5��#y��L�����
����}WI�f	Ȭ�[7��<�d-��Y5A	Tôv��BI�X����7F`Z���u�"������m�;�0P�w�����^@�#}�٧f�ה��M[yfk��/���:H����Q�VgpO���&b%!��x~Iyq?��P��K5.�xXw�bv�n�2#�G��.��͖��|��]�;�o���#^�n *�?�4�p"�o��k��}��
��{;_����9[�3��}W����@l��)3p5�3 ��L�-/��<�4��N<�yo�(�s��v�N�c�e��U�!����$�B���A�#DO��O��opa�%B����i8��g!��%�p���-+�:G)�gx;
.	���Jp��?���׶��VWv0X�k&��D�h���Tq$jj�N�*���7��%�#� �Q&���ݤ���AB��p�j���5l�Fu?e�����l!/=�Dk����Pt��{L���Ha.<B���I~+rPY`�:��m�R�vX�ad��ת	��&#�"m�Nf�Ҩ�RWA��uŻ(S��Hҽ|���[�����YyU�/�h]Q�q{������w�]���$ɪ#����I���q9���ݣ���W�WMAO@��3a�dW K`S	w���؎.��G��V��N^�P�����峧^��Ѐ��{4�w20� ��4��_�
�d�<����h����k#�E̹�,�Y�-	�*�e%ʀ���O8����aHdI�Y۞ ��Q ���IIR�H$
ɚ����¢��%��3q���;��P���$����V-%p���fyiN�<�Q`
��Ȋ�o4k�����l�W"t}�����J|�>)��Kh�I=�:N��+N��X2�.���-HD���c��F��B�K�	#ɄyyS�|H+�������}�ҵ�U�N��R�� *��w�r����u�U�F��'�H5��뚉A{c�-���R������+���8����H���JCZ|��	���@�1��N4V)���9<�=R����I��1�v=����q�
kJwF1�iu���iA��^w��J&̼��t������J���jz[���S]�A���#t�Z�d��:5�	�\Ε������ݥ�+u�)��l�'�bH�߆J/Ė	��A"�G������<d�\BH��[r\z���6��2��5�ca�8����O����p�xSK%i$��ZgV'�N<]�9"��j �wa.á��փ�D��|�a:��j;�&��
�Y)���!F֨��k�չ_�T���%�u@���F���_��˨Y޾��pp��L�T�Ma�V�T��Zqw�P��u��i2�����X�BX�B#�]���!a��V��1n��T4.8Ed�i1�91j�C�J��{3C�ϻ���~*$�^lƮ�1Fw�08��:����9v]��54u����� D��3u%`n�`�}�.s�Q}��aD�@M���h���G�7�co���I�Wݲf���,���d�i�md!]��8ڀU�h�b�j��K� �&��M�Y���t�iX��:&@�QyeNE��!�F���4��[�(,KI�g�c*��Fi Jk�Gvߗf�j���q[���[Qw�jm�'"p�%�����	���S�_��
|tM�7wI�H2N[%�I>����u���גN������ؚ��\]�௖ 0co7Ɯ+B��D��4����~�MY�2o�tDB;y��S�� �NI�
�f�d�pο�CC�]n�QB=e�M����U���C[e���9�}��mr�*9��m�}�t�0�@b������:�x��{�U�i#;P��z��-�G��E1W*����b�V�'u���0E���Kb;���`cSsu�2J6���^�#/!����h�8!k35S�p-]�ϳY�g�&߳ȧ�u��ִ��C��{Dٷ4d'̱X�QS���\�3=�&�l���މ.��ǁ�n���_\W_t��Ң�ȫ�#C�_zյqb����[��'E^*��Ӿ�����;X(?����D�vw��,�X����w�d�R����:��D}$ȸ�`ԃ��N��p�Ʉ�����q��Ū�KC�� ϏX��,�yf(�w�8̻-���&���/�ӰS����1�Fu)���;�^�B���ip�q��1��98��<}K��7��7�Jŝ�����Y&��k[�En[:%Ⳁu��G�.��P�O���c���ł�.LG���rQ�ҏ>����̭!-j�Wć]q29�\��t��9J�@�S�f����V}Yf*e��Z7(ep1d�s!=����m��G>�ѧLg�%cNr���+� �o�.�4@f���z�k�A�J��l4m��+���b`,�`#�2z�.����!�����p��x�,��Ogn��:�3g��iS��yb��ƽF���$W�	@����֫�OUzzBP����ʶ�[��A��2��l�U/˱
��y�pN�|�POѾ�Z��҈Rx���=�T�Y&>%�y���-�E�%_�VGt9K����P�6$,�F䑐��X
��;
v�K�d��/\b''�O7��Z�4��R��"��'��s��3�)R�����Y���A��9D �����H�D��6EM�G�.�k��¬�`}�+�o�n�ܶC�r��I�k;d��>�nh�q��vx4�����z��hR��.,�>	jU�υ\G�����@rSmx�b� xV�`�&n��]x�h�)<�W�/�k�B�J0�$��Q��5k9>ٲ�^X�)Q[S-�`��n�?Xec��)�H�}����[]4\�K���y,q��`��<�;&����X���zR�Fea�:&"���8�V=��V�p?�:b��l��5v|6��������ˆ�XZ�!�����)X��Q���T�䞋�ϙ�IJ�׉���8�P#��=}�`�R��sܡ����J삥��K��o^�;<���
���@��Bզk�.y��X��m�L��U�]�៾��
��F��U�?���s=�fY�L�G("E�ǐeU���uxWJ1Xf?Ǌ���נ�?)��!�UwG2��A���DU۳RIq�b0~�f�G�K�V��F�{F���
0/9&#Ʌ\`�M�iI��IaD^-_9�w��������7�~��nL1�)l#��9 h����Pi�t�~|-��y���n���V���4i�R���m����I��������T�8yʇ�~C��5K�@M
��$�:Ή�s��D�?����bJ�"�X+��Op�4-g��&H����?��䷯�p��S��#�0�Dy�%J?��ѻdQ+	�7����@&�_�x��q�W��������0�w�19+�Y��n���Oo�%�x^ȳ�Embӳ��/��R"g���pc�h�@,ʁ��䎀�4����c���1���tj��SZS9����Axj��w���DB�p��9t1<�m�݄'��\r�.M
A�4V�J�b��V�y-T^��U����͕�K1Vp����U���Z��̌�7�G���X�.!���C�<Qe�b	D2�^�-�`���&�D�:�H��.��){!r��x�J%J���M�#��3�Z���|E?wTd wX�"�Rژ͗�� �0��p�$�>t���U���x�Î�R#�R_%�&�aH�')��\�5��SNS�ۤ!��h�/�k�`����Y��F׍�����X�����;��%r��+^1_㕦�]|%��U�5�|YmjQ�
�q�K
��=�4��{1�쏒��Z�S͗L%k�!�6q���5�u�EbkC.*2'Ɍ�O�گu��d�u*���\
��`�	������Q�Ѯ��B��*0������ߌ|��9b<7�O��y����$Y?6��W���� ϖuꨲB�������>����pn����\e�W.��s� �Z�ĭ��c9��x�5�[�(ez������y�2����Y҆I1ȳaA�)�l2����pIER����$�P�U4����	��q)�.����@�o8��+f�1^p�c"!Z A�>�2�6�������
��=�y�K��Qv��Ìb��-F^'���/sb"�-d&s²k�`_)�5��X��5�	o�S59Uèv3�>��
�J�U�Q�7�lMU=��x������W�3l���l�>��O��N_�I����,�+��ZŜ���χ`����X*l.QI�)UR�KR��$+��Ÿ� |�6V�(�n���C���+1�uX�Ax�!xlFM�X�;�ͮ�< �Ә,�#<,VK����oN#��%�!�w��d�a�{�x��)x�F33͘n ���b�"�z�0jŵ��4uD� r��dcwR�.S [*�s��ӠCa�qT�{�C����ӧeІpf���X��Bʚb�+�Sl�O,8��a�/|!GǇ@e�t>n�'H��D�$#W)To؜��jI�>zA|[�h�|&M�Hm?��~�ZbnV@�{\�^EȽ��I��`�9�0��n򝲴��\Gqy�����;ͶO>�(����(�g��BR��Q�5K#��z���OT�.��#Ky��W��V#�+�3,�:>�%�����$����;�qN>�m�����t�D[\@�����_��k�����`�=�ʍ{lj8����>�d'�"�T�g��1�{,+���ޗI��_�Q���f��z�A�i�h�`+\�y��55\�s�α�ܽ$��Oa�=<�Pig���5wt��T{/E�x�Fj�&e���IS�ƽ3�5p�g(�˴�����|�.Cղ���m��^;�8�1s�;2�T>i�mt�'.Zɲ��{�m����y��J��q�BQ�E-0Vj�v2q#���Q��|��]�U�����*F�qg�J�7��e�(��w�����8܈��cM�}�x�Q�O�psH�C
<>���ZQ%�&�im��B��_q5���Q�$�gEщ~a��i����?�����yy�蘬I�Z�&?`̕��/�_���X�F%ld5���L�sʮ��0o��+MYϨ�����"Q/��7��Qs��7�vb[��;M��x��2�2��:-�anF��1�an���& �R�P��g�ڐ�<����Yyz��v��%s���T�C��\|�]W�@��7B�@�$�4d����P�!qח^���x}�t2�0h�*NɁ	;��&�o����n:`F��nD�L���CLj�ȠE���˄��I�H��b�gV�*-W�خV`�r�n�W?�H�3&�����b�;<�����k�r��M��'-����Y�f�B��[*���Y�r��m�&É��si*�+�5�tM<'�ӳ��FCs ��T�%�Խ�2^��.��"�l���L��=+�Mw`�-q"�)GW�I2��Q��/�.�������bѠ�'ZU���]�hCz\\��4�M�� ���{"9�ʎ ��\j�:m��yzU��;�5//��{y��8'g�X0��5�Zof�&-���E{��-�x��Ƭ�ij2W�v���~��l��T����	I�&�[T�_�&R��f���B�C���s����*�"�5��ԓM�ʺMR�|�6K9b����埜ޥ�-pk�����N�c�Q�cʦ#�G��{=�R���X�~�B�ʲ	2�*b�������i��tH�BT�QJ�Kmw��Y�	}��;2!|(�Y��^P�z����.�,׎��Q����2�m���L.b�������v�j~��y�E���Z�]"���!o,�����j"�)
����nޖ�S��-�;	����ʭ���pc�q��~_=Ѓ��[-v!��{[����v�+�u�Sq����ݙ�-��Y8��P`�#�'s�:߽�XǕ��xaZ]ysBMXFp����V�Z�[���	C.�W��]��<'H��9Кv��^W��UCO�HN������6�>/�`(��ȕ7D���v����D�$�X���0'�°Z��!|�\H�@tW��m�?���$mD�.���B��zh��!!T=����B��`�ßB$]qY�齃چ�;�����Ǫ�w�����k���j�+1�ٝ�I���T�н�*ˊ��Pg������'dW�b���s�ݘdn\Z`�*�"�4�G�ۀ��z8%=B�,$5.~	,�)7����@K¶�s蝜)�`I�W�������fdy'~�/��f��UQ[�O;Y�	��<�+�����SS{�@�I�8�����X;�[U	�H����}s����tf���;�ε�xϡVB��z~��"s�u��n�������ѦSH'e���B�=#�����/���RL�Vˡ���t�\��_5�e��uW���{� �)ۇ�W.�c��Wb�%]�5[��ipf��\4Ѕ.�:���2�9�q�O���-�l���C�[:��pŬ~�zB��JM,¬Z"�"�cf�͚V�Q�y�ר���T�����~�w�d���?w[@J[����MTlOGe��/��!�/'gS����Z��R�m���780�q���`��SQ@ѾEq���[T��]�UH�,q��0�&`�~��a$b��;��n ͻ�_6�	��:��Vs֌"W;8�S��A(T1������ʧ#�l������X����AB��p'��f�/}���������@NHw@�a�O�>`l�~jA���2�Ai�cֿ�Z=�>``����H���&�,�CK���wxx��f0��D��B����Ƴ��u��� �܁kxV�޾�!hig)��Re�{��@����l�cL���t��9Rk}�� ,XiL�K[q�a��q��V]0��ڗh[ڛ���X�p	I����$�=���f%����c�d�SLJ�/9x��l$�T�G�=
`g�:��:�Nd];Jű���	U�֚�����f凗�/��e=�0�9t>�����y��?�������΅��S��BCjrϣ��i��G)B~��✌����s�����	��2��j��>��Ž���%�9��^���&?�*{�w�s@�����F*�j3k����b�m=a�u#�y��p h.��`nPoDo˵�(^0v���>�xS�Zx���I��o���_
���He��%��o��@�@����^t���u3�PK�xW �Mu0��l��Ö�P�����v��R'�V.�c�9���:u!�����r�n}=2�R�c���)��h�)S�;�~Dw'L���-��K�x�F.��I�޿��g���lS\�<��7wo��d}m�+�@]PHbs<Yn;<�%O��x:�9'M�2�6ݒT���"�/�3H��(r�(~)2+�I/z'�/YB�`�]�]�<�����^Z��	zA �.9�Յ��懗��y�쪆,�Z��aA�~�iW�Lϭ�m~�#�r����,讓�qK9�ȭ�S�8o���_��xV�m�g��I3��dF��l�-��1*��=,���k'-adS_9L�����dꖾA��
��^ 9PmmWϥ�)ǩ�8
�#�u��"q�AbB$� .����vx\1lBb�v�r�0��ۗ�3�y�$��7���طl��[���rsir7�y0�0�/=��$8�:�gzjF
87S�bk�^cP���RA��@ZpVi)|菲�@=7�`f�@]��nhpol�V�XiC�ICd��x��=�"�=�
ˆo�h�~*�((�}J�����zX'�Ovla��5�p��s�u�L���Lm�%Ɉ7�{~�n���@��k�Ru�r�S���._�C�ⅻ����w8�0c��t�'��3u��(�q��.K��|e�C��cis��yٍ��~�SB:3ﾖZ�U�$���4W�8O�g"��(Y�1yُ�	F	V��i،l:����M1�O��f�~�ъ��f�X��,RT���S��b�Æy"��U�|�n�1b�˫\\�������-�BwO@���;�B���D�O���$WTQ�Tt[E��2��f���ͅR�n����Y�<���tq�K�5�E�����&��+X2V����h�T~���,�X�E�v��TV�uq��y�v���_(���v��Jɳċh�*�i �-vE��M�
�d	����MxY��|���k���4�>+|�n
(�u���OjU�E&����[X�5qZ���7uXW`O��S=��[-��(;��]�NѶ��	��9��c�`U"H�_mj���!������ɾ�$I=
��[n�F0���9�b�
�@�LvM_T�����x��ԥ�i��څ��<#"$C�Tg�"~�Xf:���&��ZZ!�7s�ΐN©�T�5Y�ϑ�9�I���P��_rk:��B�g��\.=��$�n|�SI��X�S�͓�����Jj'�S�HI�K���	.�Sa�ڠ����`�3�Z
��6�h LR�#�!Z�|s}�	k�NAP$����p��H�8�=��'�*�L�w1��F��Ci�ص�N��d9X���onnh�W�0Q�njr��hל�u{�1|N��$����*D([1AO��I��Z$`cU�8/�9\/�A��n��۸M�t��K��� ��
��I/~Zҹd��cð} y��
�߆I��S_�Or�W����K��>aQ�_dS6�KS���f�Ӟn�=��c��Ē晱ɽ����޾O�5Z^���0��<!ix(Ss`F�N�<����,͆^�1i�^�n����K[�ft����]*������4,-�D��8�z��x"�����N���Mm�CvV�b��(0�D��
�3�G��;�S=5�9\E�e�[:^A��2`�ͤ%i�V~�R����<H���(Hn�ݴ�N��ƅ32M�)q��X� �� t�Nr���ή���q����}QĞ�-��ڝ�"Bd0Tm�{!������N@u��ܗ[~�����T���͢'a�l���iP}$���}���2ƹ;Rb�Ta�8>x���#���J5}��|<��W�rm�Pf���3��u�� ,e��g٪����T��>�\/�0f�\B���K�Ӌ��BeDX���Z�Z�Ȏ%�ق�@t�@��c��p�16)�6��	�v&R�>N�ϭP��9�A �|�5Ag~���޸�E�S=7�� ]�X*�<��-5�����JiDQ��R(��y�����}7�����Q�N�7'���RPS�F��1��۽����W8f������?�9	�{t���K6��T�����)_��J���N9�~
u	�jSh���v���4�+�5 �3���3��4�wܚ��|/��@�ﲒzf�HWȐ��r0Y���02��z��A���V����#lB�ɤ.B?��mr�Y��da��0~Ȍ���)_�幵����NL���1ɝ�8��LJD¤~�n�����e�ƶ=yȩ��Ui�'������\0J�q/�3؉��XFIW��>�A��eR�)}�@��t��sބ�� �{�\�ۗL�>}�բK�
���7�@�������_9�Ǚ�B����ݹ���4ܫ�&X�)��+(�u�H@M ������?�z�Σl���9f�ԙ��=w�ᤐ����H}��"� P^�.HԦ"6)��:S�5�BB��k�I�c^[V��f�%����������������9s��V�H���X��4���k�i��Jpy����,ςN�"z�Кh��^���['xo�ھ�d�� �Ԫ<�@/G �:dBSHś e���K�k�"*Q�.J��zkp��%$	���Ŷ�DPꅭ�ll�f��+�(ܸ*=���)y�� \�ݣ�U6q;DL���׈}�?�<.�[�ٌ"Y	�h�������w��r��c&2��4�J�"�����GW��pY�ģJ3�6��8�-�<�h� �,:��ĸ���6�C��@r���G8	��m���R_�SFhh)�c�h2�(W���R�6�)�G[g�⁼�ip��ր�V��98y�9��jjij�"G�O����z�\��{#�G��㜜%��7v����8���-o+b�{j��
���S��é�^l9H#�N��5h�0��\ৠ�[]���e���ȸ�;F�p��~YO�����/b�����ۑ� I�zeT�E8��A`�6�'V��Uz��)� ��4�c��Y��?���,u��
]ME��&ш�DY�� ����<�$a�������QkRM���J���+C%�Z���B�xh��*$y܀?���[�:�]	q�ntz�EmB~O�[Dg
�*V�F���S�]���.�d'�dnae=���Rw���d��h?Yð�5D;n�:qz=Y�r�)�`������Ak��nW�XО��J��:�`k�l�9|H�|aݛ���Sgp��.G ��֤��Y,��%LP�y2t8��x�B��̺��$M���B[TM�S{ta���0��k�+zy���vp<�K�|02=�!O��4d߸�����M����e�r��0&�2��\ٺ���G�Ho6�8��g�`�����7�VZh�k�f��ןX�k�D�]��Dɋ����5�*��?��y��� #�Z�s�x-��_�{�}�[�'F�.[�4�I`A�/.yVw������3��rv%FK�ℨ� ��<�"����Z�Q{�r��rYC���h�7@�����A��&�����Hn�qTvpՇ�ҥ��_St*a�ʝg��ŉx�#(9�EI��F���ڷg��Dl�*cM_U2B��<}P����3/Ifa�YNƞ�Hp��W2�_ByWI�� �#��ś�g�M�D��.���	+�O�m���r�;�:_�"E��˕c�\����X�� �?�ј��6�ֱ��A�5,SNՇ~sD�(�r��p�9݃�,K ���ZW�qʣ���X'6Vϙ���;m��|u�@�c\��M�����:�\����A���i�`�!�+Z�q��� ��o��y�I<ɾ�:oq�\���X�^X�F�h�����?�X��8���������]�L���:тx=�{^�d,������[��4)���j‏*�C�Ӊ���LZP�d�Xb����G	Q�1u������L0:#�U����]�\-���Ā(��5��.��@6P>��9�F��Kc"k�����JY'��ѹ�v��󝪡��Q�.�Q
s4%��\�Z���S������L��xۂ昲������?���_	Ty�%��ʩ�~�3�e�W�It��[�j2؏����U�-~JO*/�Z�ɧ�p���og]A��'�4�V봿^�c��&t�^��4z��+���)#�[4�����H�T��/�@,{ɉ�D�Նa��X/Z��S�jA�(�1�l=�u
��|��3z �|�w�{� ϵ�j��]�X��J&}AL���f^�+/% c:-����d`VI�tux4�:��,��QՉ������P�ţ����7�! 0`J���͢"(�F��W5�݂�lJ���y^b�_
�(�Y?๯B��A���Eؼk�JO4�o��5�Թ��ƥ��x{'R�v�&�1�����/��KgI���U!��#��F�����U��g螡L
���Ѕ�)�}>�}�{N6,t����\��r��ەvݧ=�\Z��ʒ+��/�5?BVއ-�,�s�!�K�l���:��:6��1�B�����(��tR�sr2�4n�V�]�垯/��4���։(��}H`p�N����o-0V9�1�k��ڲ���ςyQ��p�3�)}F�@<UB���$�yT�^"A��5�=�l$��N��ɇ�������276��iOo���у3)�"�7�fbʂ�T���V��uC�NF�Sv�(/H]��d��QWÚX`�t&�B<7�~����GY�ٸ'$����t}���ƅ�b2�ŉPJ���S�6�)��m,�z��D���=���O:o�=��L�������;_��v"��ubu���y�~<S%@�E!@Ԓ�Mpnas�l;m�Y��0嶕�����xZ��c�!�C�X��zQ�;�[�-W'YP����5�~��{ o�\��]�YL;>9�3�5��f� �VݬJW�-����P��_�����j��	6uf߬z; d����y�{�E~�紊����<��[����/R�Eϕ��Y��v�Xx�i1'���ڣ�2=��16W������"��p	�ލ�ɼ�?ڱ���Y��P�~�X"o�Ͼ�>��I�����}�A�\��tuҼ�(�@��(�
(Gߒ�O����=Z�e*n����P�~D��]�#�IB��� ���٥�\Q�ˍ
x�a L��Na� ܡ���f��i�1��q�����e��[�1�}�]�4��o�(�A�XN�Z���̈́6
�^��mv:��{���I�`������
��T�"�4�$ r������@B<L�>���\�k�e�_d��l��]�"\�6�-+(Gt�q�_�LǗ����7���-^11<cusYCq$�s=1I`�]�F������&�� �q���Jh[�4�UL�j�
Nl�4���PL�]Hz� =�v.Q����> u&%����{��|�ZV����r�;�KB�lW��^�Q��@�2���U����(�w�LP�y�G9�=ԛ�51H*`UXH|8�X���6>�49��l˴���5�Fe�,� 9��Y�o�+L�A�B�� ���S>����)k�p	r�"�\5u��ah6�..�SD2eC���,�����'��V�aϥ���3�`�>x�	�Hb��$ը}�9�?��S\�(Xz!ޔ�H{��Z�e�������xR��#g���{D} ��n�](�"ui�����0�}�YI�Vdf:s�~;�bH�y�W\�Utsu(b[�t���>�N�� ��G9R6k�u��M%څ���ix|�Ѣ��a��μt�����A��Y|XaZ~em�B���w����i։0p�b��A����`��mM�4�$/Hm��>.u�rƅ��5����\�q�'����s�B�Y�0�,!4�
B�h��h����?w�1�ɀ@�=�G�ʤ^Gݜ�K�"2?�'��e������yb����y2/���`���4Lp��
z.uvOr���Z�9�^)U���S�5s��C����Yds��k���YYN�-�����';%�s]��p+-%gr��ٞ��a�8MT;��Nm�;g�������^��d��"�9;%�*4!'�¹�n���$h�N�V&SM�`;{SH[J�)��n��<{�E6)���Ht5 �\&Яe[z�S���A\͆.�$c`\�	�̎���\���I�m� ��s��Zx��R�\����\�̛W����!Ұ2��i�D��ߠ�������J<	�a�)<��c�! ��� ^w��	ٴЪ��a�������:������W�l��}�-��_i���~�V�*@p�%���e%�a⢧����f�N��T��1��������Gr��Hd*q|X-��a.w �� �U����:W�ON���N
Y��q�6M�=0�n^o��ZG�FU>�б�*�GvK�v-��5�t*jX�|k甲�����ހ �q�ǍE��@a� F
�����'��3��e��5��ؖ��FK<i�٭d�`qn�F�a��U� ����������T�K@<��]��Fȱ�%Nc�#B{����q���_dcm��O��(5��@c
s4J�(`7�N1
�k��`��cu��a��H"u[���g`ѐ���a:�縮ǰ��z}�G���pWk�Bk?FI���LV}���Z�~�EY�u#2�jM��}�0��:n��t��sʑ����T{�0���g��wsXb�!d�'��GC��ʘ����HE0�*Oe��&�m�^��r�M؛9��,�n�����9g�@=�H^n	e��(��$�H7�HJ	Cl���ֲ��fsww�W�9j�D�N�QG�6f\z�ǐ������ΰ��V��S*��]���d.����������1+�T��l��cJ��O`�@I8ڏԔ�n�G�Lp�s�r��(���e��ʐ�O�M��H(�.)�ŔX� ���a��Č��-!įօ���~=)�5�Cte%!*))��ySЃ;CMV�zE�&�X<w`upY-���b\���5<E����@���[> ��72��oH�q��c�J�����D�~�lĨ���hCC.��ha�#/����%��<���A6W(^!� a\��	�-�v΋������Bt���꿮e',y�J�	Ϧ�5,LD�0���:^��/ِ�(�{'����b�:<3p�u��=�d|���8�j��׎.E\^�N�0Zˍ��& @*��6���p��#� ^��Fu��4�����[��@t���5�3s�ݙ�g�A
|&958��~��_��2+#�j���HȔX�x�c�9�6�_?�1�P��j�E�lF����]Q�x~�ƛ�)�_�q�<"k1����Yd��*�y%Z7q|�{�A���6|���Ő
�nc,�7���xᮝF�t�n���/9�@Tz����FC��d+�ZW��c�����4{i�퓤}�/���������}T�-00�d�t͈c<�}�
7��p�œ3����:6<!��̓×������@���Cǌ,���>9Ɂ�CB�<���u<�:.�i�Yo��q��ɸ�y�p��uMM��^�/�C���-�'�[Ŏ�ҫO$����	��wg�б��0�ț����F����y@g�urQ������DL+���u��l]g"������7�'_��x���6�@�M��
gV4�#�VP���&����'�b\P±L��;.�JLԫK��پ�����1�Z{��&Y�C�)���h*����pɃ�M��)&B�1���s쇙s�t���y��6��R�e�r.����'K����P^��t�l���զ��!��1f�\��P��i����{�v�ؗ�/�H��c:K,�����x������?z_�u(�9_�M�,��h�Ds����	%9uh"�L�iѷ�8�NGފ���w"`�*�9lޫU��!cP�ܻA0ɒL���N� @�b�x�{�"�}�HҮ&T��Y�Pz��.e~��kȂK�����7�0^�w|~{\sDb1�#�+p�S ��yN��L3���Gʷ��� XzG�L�W����(O	s�Г����d������~e�l5��yP��хm��=��d���3+V~��;��(�d���Ͻ�vg�J_bs!����ȍ�����o��q3JSs%�;�q�����+:"�v�e^O��lb�/HV����}6�gb�A�
��H+��6a~���=��ډeu? Q`�L����B��D|ԗI��Dm��lH�\��������jUwR�|��W�T�&��n��Z=nԢT��z�S��ZւV��DM���ݡW.�9
���>��@F�A9��
v%�N�͈G�2�{�_����Z�fP'Z�4f(��q��ޟ`�_�
O�����h*�B8y�)�/�\�誊}�#��F����IsH�3�|��2�%l�x��mb=����z�A!`$,�W&�G҃A�����;�%d��)F o��:g�v���5 �Z���F�
�U,��7VU<�]��RU$�t���Wl�ب�+Ȧ��1��Ҫ�=���cf��z2�n���#��A�A�v�6��PEF��>�J"gؐ>�e����ƨ朄�.����A�r���P���h���h��'m���'Ν~�)�Z�dJ+5�긿��Yitu��y�o����{�vH�II�I�mW�-�������b}�>kG�	����c�B��(�QU*J�Y��Q�$ŵ��˭+���H��QL�^��ozS�췟��n���N��7�[	�ָ�����PN�`	�jkS��z8�dl�Y��ב�;D���'t�'���]'���FSP#�a��W3�;t��ɘ���Vt��܌ﴮP�#Y̋9P�'��|?��[�U�h$[�������=Ȋ��m(��W�V���gU�"Y1z���?�oh�d4��d Q/��O�h��`i��{%�iA��vS�i4s��x�I��.�@oTXVi��,��"�ۺ��F���.�.�벫$||��4��u�v�nB�\�հ���TF�_������;���Oؑ�6�}����C�G�#���>�R�7�W(��22�h�o���t��T*CY��4)��|��w�=]]�kǬ�q>s*C��bG�Q�k(
, �b�P���	K�"/��1�[�����q��b��u�����B}k
Z����B�F�Hik� {�A�AQR ,w�&gT�A�y����Gw ��4y�W1����U �ٚ6��#�Һ�'��T���b���l��k��nU�-/�S��eL��0�R���\f���Oa]��\,T�s��^� �/䟪`��;LI?�u"��������>帏uFbs����{2���[�}b���h鉡I]"f�8B��ӢA�_�&�f s��3̉6��MU�픛8+���&Փ�/�]���	.N\#�Ǭ�D���n$��TS���-۴}��n63���������͂�b�aI��g�����&u?�i�)l���JZۘ������6�Q�}����ub��4h��h�4��s��ѣ��7���FU������e�~���)��KW��aЈ)�?ؘ�[�B��U�~E4�(	�Ͻd�0�d�����n�.�������y(;�5AoG��e��:.�����p!!l~#4�w�c���m��{	�r���5��6�Q�2u�#L;?�������\�]�e���!ӷ�@�ȶpxD����������m>��(G�-��Z��3d��t��u��)�_�F0x
��{��s\)���y(9�^���o7���7���v��7-��C]��(���ֹ��"1)�Ҵ�Ur{����t�*~�u� Y�݆���f��=�bN蹿FR:�(���
2�~�Qc�t謺���Y�WG�Fm�?G�3u�"VP~
�R�D�? ;t��g5�+�{�٢4����SE�}s#ݭɤ����Q���g�˃�Q�\�����
|�#}�
]��7ӿ_�I��8+M�&��Sh%�/�(B��3���(�齾ޞ1�� �[mjM�9��-��٥�z�y�W5��/�A�ݔ��05ǆ��f<�!��MTn��>���$�>/�.'k 跛K�lǙzN��j#��!3�,��	&�u��,��R���J:����l!�9Se�jZs��a��_�Zs�.�X �2��8�p&)��?��8]۵��;�dœc��V`Ͻ{���wB�L<4s��3hV�c+��m�*�)�`I �e��2�i��q��H�Z���n����m�48�f%C>lX-�b�5�'��ۿKS[��L��_������[��'�jf;A��@�v�N�LzUx���Ӫ"�CQBѵ�iI����(j�/�(�:dP�;�װ�@Hړ�F������;��MF� : M��yA�ȸ����������̌�"K �#�W/� y�^����?�,�����I'0��6p�O���.�&yO��H��S# -��?��(-���;���0��+ī^c�⚕�ϴj�w#m���a	QG�=��9w�/�{NK[�Ƭ�����V�7����d}7���)���?>K'�Z?�j$̑�]�h��7�r��^O�aL�J�-3٣��bpFب�kJk���+% �wK��߈e����N�K�
j?�����z�Q�r7[}{Mu�Ym��!ˏUYpț �:^Hl�
��gWn+��"��Q��Y3���R��t���I��9Z�WdтVX<$���p�v�6/��wx�=�����+$x��cʝ'4�j�����`�YuZݗ3�Y�R�˰=�Fzn��޸��-�!(F�:��X��yc��B��xLU;KEĖ
�j�&��pF�� �Ӂ� �-!�J�uE��D>��Z���a��o�ƕF����B����UƧ_�G,�
\�@LT����b]P2����ެ��YN�x�Z��5��X�{��N!g���c�G�c��'�����S�C��1�@kt^u�ŭAn*�|Y��:�|� �r�V�ʟﶇ�UD���WN�nF�K�ֵ��T�_�߫�w>�]M�{?�R0=tx R����R4�$��|O��pL(��DmP㈻�q�O�}z���Y2�����?���'�Z�Z�il������<Pp.��B��Zj6�blNh-���e�	���*ש~�����痔[�-���u1⡝�Rߡ��b+?&%��mk��ާRv6/Д�#Ɂa���5y^Y�{k�V�;׼0�
˧���W�Q� �2Il}�k���N�Y�tk3��R�JUJ�T�%�0�u�o~Mаi�6�}���{��{G�m�	�q�Ӈ�O�\��y��P x>�I�����ʟ�=����i�>�YZWc"�����)v�X��["�4d�Q�$� ���f���B�s��({���f��Y�����2�A=�2?����²���Q����A��'q�8��~ֹ���q�	��H�c#rRa�k�{>����r�'���� �3p����c��S3
�lnЕ���]R��B<�Vbݣ�r�BV��P�U�6�Y쟸��Q�s��%{� )�l����6}E��r�a�}KK�!��0�-�g�P`�y��j^�k���/����^X�N*�	x�|ز��5{���ґ�se�K�J�AKy�p���L�Yor��w9fwyg��{����Q$MW���O�&���:d���Y�#��a��ȯ���2^Y��� iX������Yul��l? G���8�Vu�nL0Qud[C�Jm��Z|]hK� �3��=�ʕ�uP*J��ɴ	2��KH����S�`[�"����K�b+�D�A���xO��)S#�ܮH�t����6�?	�,�����oBᲝ��$HM���ܗ��w�Ry*�����3-�0P���T���nN�ꕬ�O��}��0e�xu�|��,s�d2tZc	����+��.� �[��z��.
\7����@Q5|Il;�����|b�G�r���C����=-��b��Z����fC��ñH��.�x�*����5�����"A�4#P��ZI���jv�#C8%h$�}�Io������u�(,�O�J}cb5�_��|��{pj�3K5��}Nﺠ@����#�����g����S�.�X�mX��> RCe*#���{7��R�-���a����es`W[{R�t�`Z����"J�ݪ�U�4ڰ��4"3;\��K0*�F�#.D�8%V1Q�{�蝆#��$�H(^:�0�4O`_/I+N�!�{W-6GB>*��k*&7b~A�����C>&EOZi�����������q&E���?Mg��HD6��g{(�����p��8Ѣ��2G�'��P�����Y��\M8幹M�f����#��#�ʒ�M�� e0a�Y�XZ.�����;7^��uM��Y���D ��"�8e3�ce��j�Hr��V�l��,-~�o)7�-dbI_�"qj�½��3���2�S?��d����sA�"s:ŭ���0W��E@^OG� �.?/S���]�6;;���,�ʏ{�>���'Z�M�B>�2���.>���'�)�Dy��Ho>�
4 $��j��D�1x2�I�-52e���u���ƾ�ܢ7�h�|��6�z]��ڋ<�s��}��3X�aP�����
�d��p"4Y�����
�y/�DCdJ�E�Vc=�Wzm ��`��f�9�A�����~��}y������4e��t0����|��h	4
�@�{��;�d���3�0�̼��>�0e_O"�0N���s놼UQ
*	���oo��3{nx�)�Tq	V�*�9n��W�4886��"3�7�,{�(��˙��]�٦��~���pH�Ѷ&I�e�P�
�7qA\f���fM�
q������J��y�Ѳ\
T�0�	&s��I�5F���ؘ cX�f��Eȟ�b��o�}�;�	���j��h�$wj^V�01���,=���&�n.�����t/Rȟ�U����`h:�Ղh��`�
�%<�0���5cda��fyt�Rj�-�Y^�{����O���}V�J��� �:k]�t�xD�h�������=+�75ʫ:�hY	Ɠ3������y[����^)�����hQ$7��5�z\!f?>ض�w���FQP3E�7}�ǀ�D�-N`�E�d�Ou�TkI���.�AMȪ;��kH腮-��|O
/�11a.E�����D}�(�nnw��0z�K���(=y�҄�5�.NO5ҥ����'�z
���U��Xt�q^������O+�^~�}t �����4�s�F�n���K��+�����X�W�tM�:ǫXOx�d�j�'��D�.>BA:F�=l�x{ �ʞ@�gvC2ض��|n� �� ���fv�ؒU:��j�₩Φ�_9�;��Սp7 y27����-2Q@��
���t����v����*���N�aT��4��PA�ޔmWkIm�L�[��b�-�y�f=��8G4���@z�+5��j*V�CA���G/Ř=�yu9;��6����Ly��8����f�M
IP���Ŏ}�W�kT�y����0�g�K�yI�l9
@�+e?.�H�0�s�b��4._>?v�W�
���ٳ
�G�D��W��7ͽ8����q?���X���Y����qh�$�5���n����OS��������Yeͮ�d�}��f�e-�O��~����{p7��X�*�����ʻ����g�ʎl�2�c��?��M �{GX;�V(	�~�Y̞(�B�'_�_TY�)st@����׻�]���_��ҹ����������5��*l|���!�W?D��G}{ym0TnEM��b+�
�q��͡\���<��4���>/Ot���-3i\�`6�r�<c
{F�!��9I�6��L�sp �c[v�u �s���/����nfZz�D�>\�ʭ@����TF��
�2�I���T ���{�f'N�Y�As�����9�<8��A��Gd���A�AH�O� l~$롍^蓷S#Snt���&ȥ v��f	X�R�"�wo�6���d�q�&�����Ry�5��W݈�A���%����~�������2Rd��Mv���	 �s���uwh�S>��B� ���3{��CR\)%cD����RDͼ 
o��2�1bp
Ғ����Ř���S{<���>��*Au��bg��ZN�P���P<}|Y�n�K�Զ�F��nҹh�bd�.�(�7����vƘa����h2��mL�b�S�wp��NF�).O5Ⱦ.!���ٴL(6�;�2G�����M
�-�59?m6>��)�d�֓����R�� �vP�l+c�P��K��g]���ܛ��f �����M�O�{9��XG1�5܉�2ϣG���[�tܶ��9�4ժ�b�k+	FL���0J�(�S�1k,���NV���\����mI�w�.a�:T0?(�	_��*�������X��T���;v�|?W;��c���J��T�d3O�����T33 ��ݎ��w�~=({���D��^�����j���-1�'��� om D,5�����Rw�H���WH��I��;J�Ɏ �f��X/�Q�1�3hI�3��D��u�=�8b� ��w�ߐe�˄�P!�yw? �Ԃ���U�j�a��������S	��R�-p�j��be�����O �'�l�x	�[o�e�/>���8��˭��m��8/�P[�I	v�ɶ���ɽJ�=i1�]�s���:�B��A�]��h���	��5������L�����Sj�����oܴ?��Z.�S+�]��$��e�:�N�H/�5���jb�m��|��,�q����	\��\)�����r����l��^a��'z	�s"�n��k��JLN�dY\�#x�|**\��*�:|�J:����8VQ8��'K3mm���<,�҄�(�(ُ�������N["'e��g�����gc,)E�jخk�TT:7��>i$���(2�����)��/\�C��¨ѢWc=��l����[G���8�ۺ���(^鐩?��;Us���p����f�\kU�d���D��/���wZ�q���||�`��ZU��qM�~a��`��W����`5km�Y��0�F�M�kQL��7�W����E��{�B�_\?%��@��o$�k薋���Ķy��x�5���M4R�~q���F�>!�W�'�
������%<(ŏ6-�5�����U~�Þ����c�Ɲd����ï��%�ueo$@P("BI� �����3_�W�W]z�}�>e�<��<;�.S��dG��y������C��l�K�~��#+]����o�Q������F���T�O�n;�:����t��c
uk��"}�?�	�Py��W�-�TnGo��h�~�����V�?>��!O.��{@����J�߯,Mw�w���v�O<<�w
�����J�y��1�����3�r�� ��#�]D�*`8�VCd���va�|���n;�`�.����	�x�%52
}X�XG��� _��2�R3 �FL��ڞ1��wx�H!��MH����s�$��g�轰$3�	ȣ�)�5H)|"������/�����3CB�����L,`M���Pf�C�;	�կ� Bzy,q��t��6������O�)�7M����v�-���w&�K��J)C.rI�>.+ t?5�� Vɚu��0/X:S�`�ܚ$�lߟ�P��βٿ"L>��r+�\�]SP�\�d1�;.plp��SC2�D1�����HY�HǓ\�R �ޢuؚߔ���R���G�~+~��㒨���]��U墣ڍX�������{xe�c_�~���M�u�|���%�*�E���� ���ԾH~�ovK�@q����jY�)��m��LWTM�C#�rf�dA`sy�L=������r/�����ڟy?0_�Uv8�*eM��_s��bK�1�:��zt�2O<�D?/��uB��%����F~�.�F?<@V�Z��h�Ȋ(�F��M(�C�B]t�7f�e�g�5���p��>�����Ц���|�kj���E�.38����c`eoH�+ت�mF��7����?6Uʦ|������i 6?�M��F����N,ò��IB���6:Uup�>��|�3�|1�\Zs���U�>sc)p�qc�?� ���]!��o]b�����������6.s$�� �b�H��>�����Lakl��?� '�A�NR>��;iBFw%��9����"�J"��U�fL�}vri�N��G�/*�Yt�V�I�v�%� ��;:�GZL���]#�v��?W	秣/y���8yy���^�#�ʿ!p�h���}\��T���.R5��~&@bhD����h��cΟ�x��;�Z󟢄�s��,:��������z;������#J�,�2ap�S��b�V�7��4�v�s|�v*|M��&��4vp�Ps�VщUV������z[j���~�����-q���}Q�H�̧�W�V+�;ޏ�"�� At��:*�Ί��b���CC�Կ�a�hS����᫒���饳Zp��ks��I���}�Ì��~9Ru�m��21�����u�y,����:���m���m�h-4� �f�L|'_nd�O#�;[�[��zH��3���A8	>G���)s�[bc��
W��ܝb�G�o�K}T���;#��D�!� � Xh@��al�W�vN�>I��g�����(�� k��:���M���X	����ɬ`lvԼO�<�_G�#?4��T�q�l~���I衶@�z��u9T��Qs�㯊Fx�=c�t S j��r"���t�Z^+����e`��ʛ8���\+�ܧ�g�+�K{'*acn*y�����;>�r�9�:-	���B��Z��_�n�E�Xb)���hV����	C^�3).�c�r��Xw�*D����AѤ��b�M5�,b�+�X��T&�����jʞ?4���N9�2}�xz_�n���{��w%7Q8;���,�ʫ���J#
q�_w���M� 7*���(���������q�r����s��l���6�~/d�5O�|]��7���s���6�;Wx������wx��^{&�lVTӡ]�Ǭj�Dr��	���E�>x� �Up�X�>��`�I|�$��6j��0N�rR���ΗM�JۯYg�[�L7ty����e����,S�5���h�E/Zr�K�M�հ��=��%��yE��ˎ�ONL�w2`c�n�e��Aa��[�Ư;x�޹��!ay�80�o�b��Q��X�殑Ux�ES���hf4,���=��\g���_l<d���᰸���Bhz����
�<__K�� %bQ�S��+����(X2���9kikEEl{2x�
O?;��c��G��c ��)�˷d�d�RQm���آ0� g�D~Qi�L\�v_���k������������]�{��t ��n���b��#$���w
����9vQչ-�L��9,d�?��=Y ID0�l�,�2���	��3��齮+ǜ`��m��u������=v���[�5V�	�æ?G��%�Una|���Y;N#��ҀEH US�:��d�@ǔ��ߡW�����.�e���D���G|v	2���_(=Q$��Q��^/��t�� ��D��S�h�셫�.V�x�Y2���?�i@�3���Ě��J�jm���w�'vA����U�ȇS�Y (i�n!��:v6�%
0'�j�>���Sd�&��B����_�@I�8�#����$RႡWvd����ejqy�j����|�
͗����>*L� ���(��3~̋7�h$%�;��q����=f�� ���a��'�^�(�X�늶�\��a������$v�>t����m��W���:Gܣ�!����;��f&���4e�ԍ-�pv�|��w5�w��������kr5+XTh���$
�mU\:���L�/�2<���I��MD��J����/�\AIA�%m��8�i�D�Љ��lv4]����-�����O�[;�hc�L��l��3��?]��8���3(v�������?��\C��C�A���5ez8��%�Q5phF����v�_M}�)�`1��k*�x|ҳ�z��yͬ�#�-M��_ �4����R��+&��? ��Z�ѵ�Y�!ʼۊ!�L��U����"("��B���E�`��WI��uX}�1�Q�ٖu�7[Uy�MT�p� �P�g3�:�^J!1��z0�pe��II��L\�%�(���n" �:W�cX�w[��@��F:������k���5�q���I#�̎��N���6���P�6$�ɩ��~R�1	���B�D�˜�
��2&cf�4�T�c����$�m�<��鄔�7g"��u�H��>y78���f���m�4	*��^(���hl�_��O�]OK�u�uǋɝ���0K�Y規�߃=�E�
X�[E�r	2� |9x�x����_8+�"fRV��<ҔI�����W��[��T�>N��4Q�#�G�4�[�s|U���qGMSv��^)���B0�p 4������rU��|�W8���jK$�=gڤf��?�+)�A6��'2$�1���=˶���*#ˏq�� ߷xU�?sN���m[A�	5�._I�^�E'�
o�`����w���H��]]*k����\V|��I1�
��񁧆��Iy�u'���DY�6B�������R%¸���R�f�>tw�G�v�>�lM��3�pj¾��_$���g@12��I��
����/"L���\g���~�i�e=��:ΝN��EQo�>�5��@!]�~.g������Xd�P���<�k$��Z���3�E:@0mp���`���-p�K��یs������{s���_��Qj��* ��[~����Y��˸տ���<��!�@O,-P?��#JmKP���A[�� o�硔��x3�.�]O��n��<E�lrUN�.�):n��d���t�E>�ˬ/��4HE��m��[����)���#AV�ⲒzUҜZ��|ٱs�f�t�3�~;��"3��NԛKx
������/�2��6@1�\����U��#hw��jצ���3�2��=��#2�A�kp�	�U���K��9l2J�a]��C�QK�}�1�H�L�s���_@P	�ެ�Pj�G,�[�~�"Π'�^�n�t����_sk#�k� �(�NI�U��S�>��͇��D��]ҁw��z��%�#����p�R��)�amz��
�F�'���TG�"_+����[��4s��/Oo\�$r!�i���;�ba��Вn�[�gz��R`i�1�{������cj���ް��0aפ	ކ>�-��T�-��C�B��̺����{�����;�g䬁u���#����!9.xa�'Y��흭�(J�L�����ךF�B���ۘ��%�S�f5�봚A�QFǿڧ��m�a�,EJ��{0�q��z�Z��39��G�󆎧"��R�nS�[1��)���jP\����C�t�*������'q��3Y;�����d/���Cݿ �ʘ�u���+�W���	q��T��1���Q�W�f�;��njfh����g�m���Vr�c�$�ra��'˒���=ţ���G�8��2��W/^̛W�ɇR^E4����)w���s��}$	e��t�K��p8k�Oď�˯H��?P�>:�v���퍄a/���"0ʠ�E}�]`[���q|e�ߨ{��t�� HRъ�|ef:��!*��k;&a<���;��שM@wܔq����f��ù��!�d�-`ɰ���R
)��+1������y�JT?��zl��v����v��� Q��4�7 bi3��rb�3� �9P�	KUWq�~7��A�O\���� �Ξ�{W����4��m��Ň���B�22R��1FC��Mk�Y���vW�o	�|=T	 �rc0��6�3ʢ0���v����跄���>��ZN��¦w>�����9��ye�	���w�ꘓ��7,4�	SP⟥'*��2�>���,?��e��7�&�";ܑh�-V����t�MfK��U���[^��*�d�f�O��<M\�F�Xި,�8Zg�&BL#���{<�IQq%N3V�X,99[>�V5-nf�G� �������sS��P;�6�5�L���#�D��1��s�A
��T�?ݡ��-|&��k���A�vėY���~6u��ig9���XI�!�����?�@H����+
�_�����.�n��+��PJr��z�@w�LM|��嘫y&�D��N� W��r��%.��Q��"S"��8��;S��7�~� .��ݶ]b�p6���6��LS�f��rf��}���&	9�ST�(^M̎�HE����J!�՚iv��`"����8Ë�ޭ�J,���#�G����B�Va�OE6�/Ăd��Kd@�!Q�Lk�L��gs�Gn��B�Q(LW'����]���m�u7��=��72�w�aԂlyk�Hmi,������0S|O��&N:�v���y�k`��ì��q���K�35�ten��֊�10"��z��>���o�*ʋDla[��F!�9󌡶+YV�1���b_2�S}�չ&Xis�I;+��b��[�����4��A�H�C&x^vK^��5˖@�l-\�=����F7�NT��{N?+�l+�;ˈ�s^i�����B'̲Y��6kd��Ņ�������E`7�����~{~�Q�?�.c�eN���N���D�N|U��cW��m
��X��b'*)M��2���սAL h��aHJ�n{n�hM�T�r�	���8���f�����[����	@�K�o�A:
o�C�ڼ����6�>�������2�H��Giv�p���l[A#�-
�$��~���`V�iqŽv�hQ�q�&���� � �f��f�Mt��]5N�V�����6p��Kl���Sd@Q�$t�FgE�./��q�2�a�3�%U!G࿝��gW�t-�?B�	�A��1�����Կh��W-�~/�bi��^Q��w� إ����Y�:/��?��ٱ�Ծ\�k�X=��Z����ZN�3��r��o���*$����=�5^�t}�7���R���x���6��֭o10�1j<K�`��1#~�7?���9���F�t��bx������}&d��Yh�P���г��
ɃND��ŝ�Z�&.y/���F�w�k�\#�ow�����:�3�v��x�/�0h:M@���#����g�'S�7�9�� �W��%���s�e���U��_�7g���,�:���j�D�_�_d��!j��S���"�]?��ڄ��q�ok��o;���A��E�n� �d�=4�!T!��ϖj>mrL���A�O���� <�`�i�Q��d��tx�xd�'>�c;+_Cl������:(�3J��q�l,�h
s�bgY��s�� ��b\Qt�=�ln�C
�T��4Tϒ����YS�w
�^�`C\��T�d�~.%����5E�߮�o1^�'A�a+p�\0I�9i�V����x�4x&�dA������K���D�T!��er#^�"M}츾K?��[�� ��Z�7	�D�d	���Chң
�?�S=�1(���v�Y���+h��1�2�.i<u�6��fMz2}m`� ZO����*o`;��	���}�A��R y[є��W]�1���䕴Uܸ}�\�'��MS�����%!�AI��a�n�M�>�`��DG�_E˝��VQ�"�k�av�RD��=7Rrm.,����'�Dh�i��� ���2�� j3�#�Xa���{�����U2�5!�>+v�s�*�md� ���lN7<�3 ��Hߟý��Ds6�n��8�J���
hy�ͮ���b�!��E3�����U�W?T~d�j����F�U>|�5��)��Q��=Qv���+i�~��h_�¼]��d1�����>�c��p���/��wCo�h��G��b-i�+<̠S�%�މ���]ga�ː�lꂷ8����Ҿ��0*��-<�^�M���LP��}(�pAd��1��-��uH#��^1B�n"�W��C:E��x��y����y��/���>���7
݁�6���c�t&���U�D�l I@��6��-�C�5 ��)}?.�e�{S�t��%[���F�>�p}�ւ:�Q0����׆�,�C�"jҘ�G��p�<��w�h2L!�x�pʯ�3啽U,���k��"Eu.�P/0�E���-�_�$(7QV����΃����*P|듞fܩ�zGѱ�|\<!PpW�O�s�ע�^^X9��bP�7��&0 ����j�����?��-"�;Nu~7�U�m��!�����C���w�͚e�*�H�&,�5?��ǀ��U�K5XP�λ�����L{��u�Ʈ@,��L�l�x���/.Y�e��a4r�#�PoD n�z�X
]T��~��k�lR��_�a�,U��J��gD8��.��I�� �{&���l�r8�"�ԓ;�@OС��|�*�׻Q�>ψ�L���΍����I���n#0#��r߫�NY�׳��� 7"�c"C��Ưr�"��v=R���g��m��hl������=e��9Fs#�#�i_�m�V��k.q�c����cK�J�����{t��R�c�$~28�z�#1w4s����ò,�'�sѠ �P�W�������*�#���p���Ej
�PO�����h)#n�����Ǽ�q��-��NH�^��Z�6k�H[(݅��y�m��&<��b��i5ɠ�z[����49�1����u��P�6��o�Z���/u��k���I�!൩��LX��~�ݜ6�JҺ�1�h$��Z��Z�����]��~��H��B�Z����~�T��<��ODl��t|K�ֽ����r&w���� �ʩ(�J�)T�.��&����G�y�S�����(�V\c}A$Q��0{Ζl[X�9�'������A:{��37'��q7�/l�$�'�z\m#���ds-��۠L�%�6wI�4���j����R+�
��a
NM��Y�%��mr$y�؎k���4r�c�2���G�Sl`���۰BZ�QD�!�=|�o�8�-Fp��d���F��2��_ �hDK���r��n6��X	�����T�7�*�87(����M�]���% �;,$��5e�̗�]\!�yh��"��M]n��|��A��.R���Zl팸�R��hJ��"i+�����)����-��C*%g�JߍL�q�eܾ r˿�dF��:���'J|�P��Z����u�K�����e�G�M��ͯ�'�V�#�P;�H�}z^	�G/����W*/��TЌ�h�����v��	t�ׂŴ�m�����N�0�*��oӼT��/M�	�x��wl?��'tTrO XΏ�Ն,��k
�v�? {���*��F��y��[P܍5�ؠ���e���p5sхxӸ;�sK��I�^
D-�{�<�}uO�	�+P�Hp;_�\j���gV5��������Gos�
������VKO�鉈��GDBΖNs��*)�c\�(�,_(BD8�����Г���콟i N����/���b�B��_���rPyDw�Xkǃ(�u����
<tЪXJ-#� �f
K�v�_!��Q���@���Nk ER���%O��!P\fDq(В����<�[3�q���%�(�p��f��eEc~A���F��˺jQ��̭g���Px�Лz�O��`3�������x+ʽ�J��$>�����[c'��#,���{6�U6���u��}Fԛ4!�����{��Q���E�)�PCל�]����U�:���ҁd=�Aߩ���\��k�A9Ȍ[�
/kkdPZ�iϊ�l9٦IK�h�1A)�̥egբ��fgnҸbv7�:ۙ��*���!ތJţ�����u7��`0�.�1G�^`p�˸rE{�,���2�E�3Ip_���k������%�g!��5� �s��'Ȣ,�qq/$���m���2@�����λVrz�#�_��l��"d����mP����H;HJ��z�q��J����/m�Ѿfuv�ZQW�v��������N2sT�t���Y=����4���a��T�b{�8�	_h�/�K�v8��ōr�7x����Z��se㽨���w8��~J� gߺ�.$m-*���<�e�eo�ү	��~P�Z"!��+������{f�T��"�aݛ]��B��R���z:�y���N'�G-^�r{�E��x	�8�x.P��5� u�~	��y��3�F ��+��ڣ��@���M�������x���ƒ�����4V��e[�`�K<��B���`��wW��w<=��~����w��e�8P$���p7��� ķ������yNwFkb\�^R��xA�����8]�������)ѳ2��;�I��;����!Qh�����llvZ}f)���@���jS1�<P�P�h�]7`�-ĕ��=x
���ȍ�!��9u�� &�2A�N�!�%eZI(�QCrW���p�w�=���{s <����Ɉ��x4�|m-@t32�d�B�'��$�^�I�5�����-�	��0�R���j6I��r�sf�VVY����=>�Y�#�N�st콗ʋM���l*?1��_�t/:+�T"n�|.�I�N�?�C��_�.1F">���Ɔh��*w�
�̽��	γOFV)�
(��L˯��J���{9���8�+z�Y���ʿ"�bRE�����E+U��8��C�&���k�c"t�'��^��1)Sʨ�+�~�� ̀����_��@9��U���{�_��/�����&	Mո������~�������P���q�$���jX^n���y%������>۫�<�喈J�S�ۛHX|{�/4��4���q-�'65BG�֠��zd?����%t�BK|�	q�υ�R�1��	-�� �Nf�α�G��s�j��/_���\vC2�%�x�'��
G�pVFRd8��޼�_<Ɔx��@�b�!�&Bf����9l���]aѽj�~=�}����I���f0�~E6:enH��=�	�!؜I�TV�x�?�k�+�;�LHm�Kr�x�Ǌ�*,�Ue���t����~[T����*hp$<��G�$N+Z.�
��P2
"���B��V�4\g��ᨂU��3u<�����ak,� .������"KQ�AJ� SBMZ�����z�(O����Tu�3�TZ� �(:�~�b��H��E"��c�p;{_�h����h^fy@.8��v&&)+6b�D�r� �%������$��vL~���@Ծ�཭y��lY�j�]L�96=������?�C�9������U�I\E�K9���I�HV�&,e�Ar��%;�[��ow�O��3��]x�s.��:;��l�=��xD@�;��E����&���Ɇ>2�RҙK��xJ���[i+k�ۉ�c��O�*���"���b&"�m�sƀS�K�0�7`�H_N��4Yq6Zd5/�1T�����s�i��"����o��HnD�]��a�����MdNW*)��Mn�I�l��9�c� �5B=�Fr�^��;9��\f}Dη���11�j�_m����H|�޼�Z�&es�+�������/�O"�:A��)��O��U����V��sU��~�i�r���������9�7�)����(�ko�Y۲k�7���Xu�ʮ�Gro�"�-/���̖����g6�V�Lˏ�7���/�x���ATq�pt2�P ��=�OoB �ݑ���X��#��>k�����2z�,w��.u�q���7�%�!F6�i>�P�r0@@��;��)Py�B�壼h*�;dJkm�)ÐS��ICj6"��*�:OU��zP�`/W:2V���>���B4r&���_�w*K;�Y�g�::�}յmx/dկ�����I<:h�n��Dɒ6�z��}�X;����qäk#�@y&�w�z�}�:rP��. {���%0?�<)Ҧ�K����@�KpV�<�/�M�~��������%�R��ي�7F/��#�ٍ�C���9���N�D��^q;q,T�`��;�D=�p��IW�Z�M����m�\-'cБgؑh���I��Q��&[]Ib'z���3ڡ�������+i�f"W ��R�C�B<E��o0�9)����.]Z��M/�9[�A�e��r�~�%D�;Z�&s�Hcי'�V����&2��Q����PNGCy����Kjr�O��'9�<�ߧB��v/�n`��z)hj��a��H��OlYt������1��-`;��m��p�R�K�PN��S��9�e�Y��Ӑ��=A��.}L�'�Y�c��s�5t�bw�(4	.���XIx&�|W\{���4�+��^��R�9̮J� T��b��rN`ab�^Y�&�r���A��[�V����q�WЋq�g*(	̉��^+,�5��E
+s�gpT�a�_�.�J�j��d@Ƶ�9?#���󮹲����:��U�W�
U?��JhWW�������Y�U�xC]^�<6iI1W����Q��c�BL��3�'��	�#�����l��˙Zq�~�vyf�����B��K1�I�eU�w�6�z�z�b�y�X0\�)��]i���W� ���k�o��hQp��ǡ���aG,�ݏ=}��G���I: �������;�[�$^Ӫ���|�i��P�'"@-̮�t�����#J�^���|#Qh�"����Q<a�ӝ�D˙`]��N�ݯ���U4	Q��B$Y��J
,�J����7cJ\�m���컽/N�����,��ܫ�%�~��K_b����D	!�:0`2jsl���h���E�W��6s"�~�@�=|%ҵt�ykC.v��������_��@Q[�k��q�b�~=j	�c�~ER�k�у�Y����Z����	�~z�Ftږ�s�d��5W�


t�?gũ-�d}{�!��o�=��|��7Կ���x��l���i�����z�^��7���H���m<�qே�pS+�-�\(I(w�������W#dK�s;�u��s��f��1�D�#&���MO�'�S$�g��[�N�]溇 ���箺d�1U�?w������Fx/��;�s����⊕i�V��F6�ֿ߸��3����V��a@�;l�S��	݉�UN��&ISx]�!��,��W@�>�S�p5�ф���T�'Vnd�E�:#NC���K�������L���\sTx���Ph�����$d�ر��E8���e���+D��J{J�񧔣�����i��:DВ~���i���Wc���	�	��u�_�!�hJ؟�!� m7�����͖`�I� ��.p�Z����審�j�Y��\����z�`
�.����E�@�e5]9�;�з.^v��7�|Y����Q�]��ɇO�s�j�����"S��&��	�+^��qbZI��Rx�Qں'{��|{�ߤw)F.�U�!SR�[=Y��E�o�6��c�4\�EE4Gz��׾͝Ҏ�y���Xu�>��}.)"��d�j���q҈?yTV��K�:�ؕ o����
	{�x��������o�Ϋ�=�tK4,�0�4Y�&�md�I��FtC�_&=��o{oK�������[�����mV����K�|ߦ�	M�J�ro�I�S}��B���Z�*���M�/�V:�uIt�A��Q�=�h?uԚ��Q�3�s�ǜ,ب�c��k|�xT~﫰E����e�S�4m6�іp��m�~i�k��n'����bC�èZi��1����`%�+�������&Kb��d��ѤdĬ�{� �RRޟ�;!Ti���m�;�`����n�8����4��ۇՋ����ԥ�@�b��݊i��G���ƣ����!��7Y���&Ɩ[y_ki�nFp����抝O��`��{���9�x�v����Řϐ0b\�M��ϰ�Qq?�^.��d�ho-��{�{)�K`ݭ��q�6��2��P�~�
k�%Ԝ'x*�?�'�H���f�9A�?`����i�x�ҿ	��
����?���!Q?���h�yqWX�zo��EU�qݤU�/lk]מl������J���j��#ks�(�_��j8}�7�~�W���I%�ƥ�>���̑Y2A�fl�=����{��0`�Z�U�͖*��Ĭ�-�,�jԦ�o�[1�E��S)v�^�?�'`�(�#*D�����Ϗ_a�Z|T?QjlK��v>���w!���g2�M,��x��@!7=����[U��%���;��{� �ҭ�<�_5^Lsj2�s-D�耙p�İ"���gl���uyD��
�[:]����uԫ��N�]]��2k���0��S<�f� ��~�;[6�"�>��4z��yBӷ��܉I�Hm}_��s:��1��*�o�1�~X�<�`�� ��T���=>�X	�BB���}cRu�`�
x�I�>{�jϯ��Ԁe��1wJ2��xQ]��m��?�Ą�jJEϧ�H�:�l���K��ί!����g�6�6Y��ҌE͕��w罚N=�\щ��1��&W�w�*�6�VG ���,���i��^Z�:��0�饉TnV�%.��.��M����Y�^~n�^D���c>B��ǥ��v��&�z�~S�,^�ZӀ�v�@R�Ų�_X�Y��Y�P��r������E�րl	Q��c���,��� �I�pzbls�R��3��KWE�
����0�}�bN�  vq/�DZ�UV�;�5�i?cW��#M��Ez�����Av�\��&�<e�F�)��tA���F����
�u�&�Ne}���jF$v@-<i\���,w��u@�͒<%^����㓬)0%^D�-�N���8�	�F+��oȪ�L-1���C��'#^KR��E��0 �TΗ���-U�E�
��b�g(�^d�J��^\9���9=�=���
kJ+�n�NP����7�]�-�G�8&˥6�z-%^|S��|�J��
N`�I��m��e��ϒ�ܥ��ޅ��bzqI�}���Ĕ�:D]�+*�����!}(=m���6X��AK)�\�'ފ�j��C['mڻ�$���Ҋ�Q�7G"����H��-%v��:���%y갽��IS���3��^n�'T�:e�j8t�=��)h�a���E�f�ٱ��X�B7�O(G�6�@������]"�5�O��Ac�J^�D���ʻޏ.��z�мhґ�#�������9�]K_m�C��@��R�^��[\o��$"Ɛ{�qR1�c�n�^�D�2�ܱ\����;�;%0}d�XmT�_�jZ��L���A�����R�c1�%��d��A��鲕#�Z�Z��MV�VϚ��C�`!-2ߵ;���� J���r	����	@s������֡��л�g�(WG�bc�8͌Ct[�&.W�'�6Éu}nS��L���=�L����n�v�$X	X�BqYk�R��:b:�⎩M�
��:��}������jq��>�F��ځ�nԏ��y���Vd�4 N�u>��3�gt-f�zD��T�����!�0
�l��D��U[�A�i3u��N�L-����F��Namh���~P�����a���殸d���J� q �Q�����ȿ�+�2�9���fl��_4�(���]!�����T~-�O Rq�_CB�K^��}	�� llBtS"2�ӊJJ:��so��s��0���9;��_�bڹի�q X������Jv����84I�����CY�Rn-L�]��r
�uG� ����}��UE������1�����i���Z��u����z��}��Ȱ���3j�	��
�c$Ls)�����c̑�~ȱ���
��Uw�`���m����'hu��7>��$�X���3�lGX�N�N�й/��~h#i�����&I�ڷ����r%�����7���>*C��1x���ڰ-Z��/bg�ڪ�	]��id/9p����(D3�(�m���^��f����|�Ϊ��r��	�{�W^�ݦ�KZe���R�jU.ۿV�u2�	+��4y��e�AY	[����)�$�RT����F �G[�p�
��J��3Yyj��FX8��(ea";\���#��#�!�-�mm���+I�q��8���%����lA�Kl^�ǣ��y�P����h��ay�?���I���4�(��-��|�W�1L��GZ�+��li��������"�5���_{���݀ۦ��ye�w_Pխ{�:�_a�^)hxe�%uP_b�K�4K@����U���`!��3��}�����D���}�,�1����["�,/3X:�m��+�f���?��������F$����y(�k�=��\�E{���=�[ٰ�r�ܝĽW��-�b]��^�aY��\&`._>]][�OȨ-7���R�U�CRL�Zf�c�V��i9�q�;��\�5�`��DZ��"]Ts��eb��O����5r6�`������:_
!}��"�t��G{9YuW'O�&��X�ە`�Q�\r�-77ƾ�S�Ԫn�hZ���O,�<�Ve�� �����l��;ޅ,�·����o�/=/�%AN����{U}����>,��m�͌����X�d3�a���7`�k�(n,�_(���v�쏘����4��!AQo�`ܞ�'��������z;�/�X@TX0t�r�0F�w�ڏ�&E��s���Kr ��>ͱ�p��_����c�$v��{����<����1#^���ˑ�r}��mvAY�?�Z^��ސ����fj�y]�W�|x5�+��O\���W&�%�XM���cڔ��V�z���e}� mp_�K�ޖ�'���U�z�<�&?Y���9���t��2Y�*M#}G����p���#ƴ�+"����?�|�78���N�$�Pj��fЭm����*�`��ٮ��%�D�-��^%��0(ms^�+FK�L��(�9Dg�	}n�<;��22 	s��d�?dJ�t���Ԩ�4(�W�(s��B�I�h*�I�;���ks��i��v+�3�4�c��[��F�_d L�XҕS6�Aj�R�;� p�B�6�hj�}�}�#*rx}�S�ǟ��P��\{|^�w[)���G��/rw��P��I
���-���{3E������S�n����dXI1��`��p���N�q�qn�)�lṤebow�v���ȴ�
t=X*��"�������?	�f+�P��G��;��0�Qd����ZX���vlΠ�t��V���V�ƞ�"�_}%���#�y����$��2�k��p"T�iu@�#�ڼ����zs�V%�.�C�N�T~�Y.��<�������Cͯ�ǀ��B�c�M}K���}���\�?���i�O�q
��Ƽ��TQn�ӓЬ5�!�
�Xzv�e�;m��!d�
�7"�
G���G�咹/�)�� ����շ�dy�K���ES�	�Jm�c�H�ƭ}^W~����p`z�� ����U��ʼ���-|�X�����Z�0��_�
�q��ޠ�y(�=�֕��d�BF�Tѡ��Bp���z$�C�RU�TQ�" (�V�"�/�Of�Gk���`E��AD�:X��X�J�9i|e��D�a�i�o�'bA�S�t�r56�����X/�G���RZ�ބ�`(3Q�?��s���U[���#P,�
�l2�'AU<��cl�`'� j�=/hU8���!\w*��\���D�R�;*q� b!=�>.�1X~�Ni4f^l �fj����4�I�*D2D�}��x+ɒ���%F��D��ˬ��Q
���Q�<�b�H�"���"�A-�,������8���uyP6�5��4�=]��C�D�J��:��B�)�6��h�8�΁�	�`���2�f<��>Y �7d+jc&N�,i�r�'�Ӝa,����?�J	WԄN�oN�U��Kx��+��|�t�a��Vk�,@�v%��q�F/���r��!3� �1�~[��Jz�O�����"s�Z�A)����X�؂�Ӌ���O����v�M>���c1q�w?aً( ڗ�J) �z �YB�Ϳ#��F�_��A�D�?�V��*ۮ�Y��t�60�2$�t��:���?.���B����<kN8��]M��������RPz��T�ax�/�)~�f|�A�v��FH�'AR���\�Tî����rT�ى\QJ�w���8��:/c�M��6?=o�T*B�S7�^#���;�{D�p���z����>�K�<6����w`L�h(�jO�7���8Y޼�#���u-)/�l��?���}]�=�z	�Ү�}@/"՘��j�^��:�!�N�%;�  � �ǵ�KAD������\�
��C�-�������y�9�q��,�����r:����-)�N��X�h���Ѧ��.AG��z��%G���aZ�lm����	���U�X�8�Lڧ^N�1����� Q�v�ATzJ�!$7;�ڳ���3$�YW��i|`"}�$�0�\_��e���c0�#6����mY�&�M0���T��-�+�TA�`����|0P)�����8$��`���@�M*�E��x�AO��/��0�3���U���D^�H�j�e�jۈ,�ų��4VS���(6=0Y�O�&/�����,~+Y'$���eN&�	<P^��vD�LD�t�܍N&f��I��t���eyl+��q@�N� RS�m�Dګ�\3����;�R�(�s߀��)�5k���&�v9��-�M���i�Jt���?</������
�@0V��L��o>�5��r�Ev� �ȉ"��׃:-��k�U���o������R7Ȉ�[n*�o#�p	C��6��0�8�<�C,�q�<����	�"2I�.���d�	V��3���l��>0^���xD4��(��pd�F{ӵ=��=���{;]ݴ���빰�_]������יߩ��VF��^^\�[>�:n��ua�cЪ�R6�Ux���$�����gC:~��Wɰ/�8��sn���@����)`Ͳ����Z)���]�|�"$���^��i�C#�7#i��6������s�~��Ҹ5���~5Z�)�t�c#��X�$r�Ŵ��@ן_�b�|:��PaLE%ƊO��@~*(�=�ID <ȍ�)�+��Q	0��Jm+v��(�Qe�E>U-H`���WH��Y	�3�g�~L�3��1��f̊/� d�g��5��S8��܅d��ooW;0<e��NxY�W�t}�OvSk�زŌ�����@����m2����v"��E�-�W�e��``�47�S��Xߙu�d`��\�������!�ػ@2!���ߧ�k4��EA�K(CE$r%�����gS~ҧѓ�[���Q۶Wj��˾��OWhy�lv>��r��\<�O�f�pӀ��M�N�T8�-��r�E(^����9���{��n�k�0���Y��d�d$��WrY���%A�5���g���e6f��|�0��S>��Y?�>�iI$r5�@ve+�&��J*8p�m��}�5 �w��=�z��?J�Z���q֠��4AJϮ���%J]�)�>Ο�~���օ�`�;��/�����X$0a�c"�c(-x�Qz�,��^��5���ٌ8��a���U�3n���D���Կ���A$pMA��luP���\��:���%c���|�����n��K��JZ�_6Y�$+ʖ>��6���`�H��f�(%1����6�䴯��?�C�s�P)��(�����<����X����[��-e= ;��c'�N0�Zp50���d��C`��T,VQ�`}��&#����֡Z:qh>�R�>B�G�������KL�P7��ۣ�B-�v8~�>�n6�{�m�q]_du�$ۣ�A l�c��CG���������xݚ7�PRH�3��B����3]Zm�"J@��Z�̧N�ɏ���:0��6ںz�^���+��_1N��8ɟ�\���}@����h3�x��m�2��'b�K@`��f�J��[v�*��V��
����{���([a3�hB�yRf"r�ln�a�2�0�jx�P��9�FZx�qL����w�)�@6$��wLA#��&SE�⽬K3� �?T�ˮr�Ƞ���(B{~�q���O���>:98w�����<���X:��c�������T����f?u��b}G{w�gH�Y���ޓW�U
c#�I���'ӅߝN�lҢ.��U2��DV�P�}�ID��-�^?�w�@ܖ�=��7��-/���n�%gH,ӿh��&��T_(��լn�C���k<�cn���;���T�R�m=v��m2N���0Z�w=�tR�;����I�mR��[��P��3T�����5��k�|A�
�LE� ��iQ�1�ޓ��aF�<����(0�$
���[�etKJ0��''Z�`��,jۘ|�E��#\p����E���C�C6v����r���E&>o�u�n����}q��05|���;}�¶t[���t!p���]F`�B��K}���ː_�s�(�Hi9�f��^�~S[6��ЮX?�oZ��z$��� �Ƞ�H�����t:y��&`�h����N��ͤ��)g�N�{mK��A�+��Q7PW�;D��U*�������ڢ�h�z���<m	����k�6ɣ�|J?�Hn�SQ7��h��P�}UY�����헀e0i�$�ODGqg�����%L��صY4�<��g'S�l�����[�r� a^Y���K|KKm�V��A����9�>�>��z{��A��6���wY��>�S|��/f��h�5�x�[�����v�y
��R�PUv%vX�oA�IÔv�XG���$bP�D�dWH�{�C�K6Pjr�JÃܫd�Gt5�O)[��6����o ����d'w���2�	I��T��z��.-���&�1+C��a}(w�������t9P�����T��@ފ ����p&��ޔp����}���u�*�U�C��?�eV�2�-:0$Ȭ�h����p�;:^�C-��������Ȧ����,�4�{��B�'A�%Y\�i�jy7]}�x�Rj������,o��⓫:�Q{��v$�y���e������ ?��(�+\�A��f1�.z��$��%t*��f�d1�㋗�jɎ�	7�H��9�{�j!���C� qW��۰�Ɵi�P}8�aL'�Od|jJ�r�mAjqi���F�0ڎt�V*�L�v�Ǒ4���Yy�t�%�[V�Tۈ�K��#&`��RN���9�˚?�����*ĺ�1_WW#�H�~���g��o�J�R��+m��+�&t�A�Ci{`w������b��/�����D���4f�o��
���f��_.��7������Ag酒Y �eE�4?/�텏��K��+n��!�P�X��B��I]=0"؂��{�s��ƴ�޶�ERjF#X5�^�e��'-*E,<	i�I}Hx��8�F�*�4<-"�	���n6�_�`֝}6��i�d�Cl�9GV��zr�Y]uH���H=y�>s^(�|y��Y��^V���Q��H�8Ȃ����_yZ죇���/���3�Ǔ3�W����{��|��쵩D���	�|�d����j��VѸ^�@�l��le�+��x2� e��@~����(����]�=p�v�@c^��X�h&K�D����:��\�8p�1	EaU9 +����h����#Q0���b[�J��x��%�>;�+�_~gZګ�������њ*)�N��u�kjwѹ�Ģг�²(N�����]i+OI�!�f	Ѵ��1�eZb aF<�r/��ʑg#�~	�3��'�Ŕ�+��*Q�Ԇ;�uŃ�L���+�'=�����M1�����*l*$b�S�3�Thy�w�o�_����M�\���;��Y˙]ם�9��Ice;�UyR��4I���������[�D�u�?��#��m� �8��Ϲ
�Ma2v%�a���⣅�`������݄�uCG9��^� M2&]��f�'l���4*G�Hv������J�k$����w�A�����fD|7.��(�Gq8Eʱ8���mm�y�b?���Oc,a����A�i�a���:�F��"���/X���=� ��(O�\��*7^*3�@}���������z��5��-%ҥ�ee3QA^�W,Zv��,z�0��{ʷ�LMJQz�N ��V�{�7���di��l'�u@�jƇ���.���]n������w�`ݡs ��Љ���n�;��T�`˵��XR��#�(�";}������:�������G���Ԧ�<�it��I��69b����l����{�~Y.�������[�"��[Tk��ZY}�A5�MJ�&VQ�.W*��p�ם��\jo�!伣� � 鱻�"�%]M5�N�ũ$�| ��ҡ�����D09�	)uz��h!��.x���<��R�����2��N�sȆ #��������W��#/1���\A�9Q�og�Y/z����z�`���!)	��� ��0��Ex�ה2��.��N-�SU*?'����~�¯w�g�D��U]J�g/�P��GJ�d�b3��7M���:?8��m�T��}p����<�2�%��#3�tKu����z��� p[2��У���E�N��Jv��>�i44�ύ�p��zN�]��B�c�`����]�RJRa�W�e^��:���kn�=K�f�E���g��B�ƪ�:j�u�]��`�<L'i�ǰ��N�J0iR�~�21Լ�޵���v	�a(̿IɊ5�O�U�I AUT�rz�@��Q��F�R�P��#b�D��AP�+�����X3�N�9�s���?�:L�!b��s[�'��n>��'9[|u�8��Nw�/8���bv��}Wc}F�p�l~Ν��-J�ZaOt�.'p�=��|���2��F�� ��3f��9.�1��Q$�KO0�-�4}_,Z9$�������r%�{g*dEg/2��u`�c�#��q�^�D�/�s�������fdY���_2�]��{b�4�Y��?�h�:qF�7�Ϙ�b����	6���P�T!8Xyf��tl�d�Q�6�����b���~�Kp�޷,S��f�`�G a����>R���lz:���Ŧ���p��Q�E�{<�u���.2��s�8�o�#�z��� XBu��3g�=@+MW�F�f�P%�H�V�E�|�m!�ͥ��@w�$��Q��/���J�� �1�������t2z��(0|��T!�J�J��`�9�Ti5��� bQa5�8��&@�]`�<cŶP���;�V���P3�oZ"��ǽ:��6�������F<�%�7�<�F咏���vբI�jk�?�x��������%C���c���+�w�x2{�������iD���*�*�[�*���4D����M�� ����E!A|7lf��O����8|)��m����^4���/�d.D���@�"�â����_8d��P+<b��l��9i��{�<#xc��B�#��&��0�܁�ԝ
�Ħk~8�}�6f��� �vd���Gb�,m�����C��/�ʃ[Y���y�28���F�!�2@m�K1,�������}9�(��m-d2ב�{�:{\�Gt�ϺLL����*�����,,a�s`!<c�ƧZ��Ђ.� ۵8w�����}J�	a�t�C�����1a�1s* L`�������8յ^�]��z��|�mO�G`�[N$$=�߫vt]7��^vq������?�o3^�f� /�q9�5Z
R隊��d�Gғ���#C�A�Ϊ�8�@N�%�t�m��<}u{ˌ��7Q��3ʞ���@�q	�^���@'�|[��2q�`��j/>b�?*�� X?���*�h9�̇SE���o�]�dz�ψ{��!�z�v�Cö����b��4�ΧZ�g���j6!���@f�s�"�B���v@�	ؕ�˴Y3�t;��2H�@�2(w�EUY�,��66dZ��L���t�S86������<ע�5<�FT4�����]!���ʠ��qP�hU�9��4�kQ�&�o�A�A�132��=�(��Y���2S͔��?�!XI���p�!�@�������_$gZ�K��u�7s�6w8}��)
C�Z������V]�_	x�;�\g�x��)V��$9;?�Y�"Ʊr�����o2�R��)l��%+ǴCm%H���D��+�c�b�C�0e�L��HKE��ݳ��!�(�2�ؚc�I��
0l�AЕY�͍��ׅ4(OE�x��B�j3p@���_w�7_G[���m��)|�Qu�Io!�v�+�P�
cE���B?��'ײ�C4Sw-Kɛ*��s&T�PU6�P1�:�k�}T@2NH2 ,5��&U�S��:
�T���^Pa�].tJ|P��k�DT�nZ��X�w]�_ϴ����"c~9�KQ�>2� ��U��m�v��A����&@�$4hV�-�$�9� D@��0M�M��x�������q�p�񰆚��t�i�a�3J_<���x���9�a�����?[�g��d�D�
�X��ӑ$��U�0%�C���G�v�P�5Tf�a
4N�����
�0�j�햌O��K���J3�
-<�f��`=��7ekP���t�ŧ�'6k��)�`��V\�3���W�����(D�U,�W�H��	��"��Z�r���J����Y!05�½�����-8�$��)~_��ݵ���v����<Z��7�]b��](��bŔ�v�^"���C��xr���XP�,>R�Z?$N�R�ϿYH�s��>�T^pE���l�#�2�x?4<�L�'�VK����L��I���[�wF2�'��7
�3��^�Z�Z�J���y��dp���B������c]q�H|���'�ͼݔ�X09�	�ç�ū��y/"[_��� o��=��+����J��)w.Pr�y��M����B���y)8�KC5���M6��q���aR� �C��߆�/R?�A@�D2�
�G,���1K����ӆ6Kh��yɹ/�ѵFyg.����yL�Ĩ����8�;�:"��� � s0��KS�:�0\���X�=|D�@+�_�y0 ���0�?U$~��m��	7C9�h���M]�[:�xN#��_�nMT2^ڏ冟o� z��R��B�AH �7�rEڅA41 �_�Ȼ����ȗ�\A{�˱���xyۚ��Q2ڸ����d���l=���YBXې�ٻO�qI[2`��S[8e����^��h[<CCh����h�Q9=Ւ���PoL�;���?�fG�h��N�k�n�PM�hQ7��b.�$��v�� "7M4�?�h���if����	�!��M�6C�5�<q��q��N=�l/�ձ�+��.񖿏sjs��7�^�G|����w�4�3=��Jr|ei�ym������� [N��
�n�K����T���W\���v��I���_z����B��u�[���s���8SP���J��sV>�IT�!�\m�N�E�_���|����%�m��i�e������O\I.�#�z��C���n��s�$��.��1yn�J����*̿�C�I-@:�j6�,^()8����C9SR��g	3�><5d��)9�9�i�����ne������w&��M*�]�i0��BD8RHP���7�JSZ�,����x�M����b�Ny�T�v����k�-���r*-<'*}� zÐ��]W�k�)��͞�h@�n�Cq���,�p������ ��:�%k�?�j΁(��*H��h�թ�������$�v(�X��s�'��@�#=4,�ZU6~����%�5%e��O-���J�6�=�/0�a�̸��P�$~����ց���F�(��IC#���=��o�y&G#�?�!�i�р,���QF����ͦ��b�*�����ul��+0��# ��m�מ]0�]�L5�}����wY5Ǚ���5\�P��ب�f�:� ��B��N��'��L��N�
g�O:�gj9�,Պ�dte���Gw�y�]5���'�X)������i��#�>���j�Z^��cc���!���C�ɎR�:��ex@���l����t�:����~LђAbC7 ����S���C��jjj�i�u��0���ZV�!P� ��o���� �} c��vJ<�"ڤ���H���ڹ�"�*j�,�]�Yqb�؍��Ra��x����n�R��V��UwHv���'U@Q�`,W�R����	<*�O���ׅ��K ��*a��-15Pj��$���]�$�*
<E�؇�̳��0A_�7HJ���OJ܏e�by���/���$ш��!o/\��F���,<�n��%'�.)��e#�����x)"��YUۀh��:��f����Ypݱ����q��7l�$F���F���L��zG +, xڧ�7[>䇍$�\�H5NG�3?t���[`(��*�|�?@0���urX��SpB�t����2>VPjz��c&�T�c8�p�.�3�`{&z��	g���{Ȓ���,$�ռ\��o)��ũ|+�ty�(.�5�#�$����0V��5�����1���pl��g& ��s-�X'��m ���T|Y�/HP�'��J|������EJ�6D�C���B�A���>�7�2�m�X쌥Ѣ����(�x�t�R]��o3\��ĥi�8�9O����_2~����gg�u�L[,��q��?�O�sݴS5��(a=ע�\���K٦�F�__&z�dU��w���S���I7%N6�|t@����n\jRp�4n�]����?���oXѓd����#����B:nf;�����}'\c@c�T+�L����<O�V�{C3j�r������Y�uZq���߼gA<\.��s�|�T�:�i:ڰ�c0��y�m���=�s�|&Cv�(���!V�x���jĲ��
�Z8�*�^)6$���,!�<�����)����w�(V~�:v�����ųR�]v���*pz���N~���I�&��o��j}�(��r��p�ί5�Lti)"���!�*}��v�n�bȣf8b��O�D�B��5Z�����^;g���K��%+��x6����;t:|�6��\�����U,��S�B>ݼA
M�B�SO��L�`���t�e��`�u�L6W����J����ϕu��R��OC\6@V6MO�B7C�lCߥ���]&=��A�(�̦R��*�g��Ļw��q��fK��>dvU��0����g��T�K�b`
�D�!��$�����H�H�ֿ�w:B��g��.��6F/C��d��x{�Wy������Ŗ��(6U�#Ѩ7����I#CP�4�1��$�S�j�Y�A�y���?@��oc�5$���b�,f7[
�a��(��d�ku2��%���Hf��w�_G�"Nl-�;n��vo�gDR�D����2�"�R�\�.b'KB����4-$�(U�b�����@�dřV�p�xf�ۀ�����¾j��Ey��9���P؅������䏣�Y:6�)gE/�ĭ��zg��T��P�!��{k|d�/,���ޮf���p�l�}� m�@:T���é��E/k�`�r�92M6
����J�noZE�S㈍�����ʵ;{9���L�G�Rbs�{N��ޢp涊��+�	>�D_0Q���9>�����F�f�����KV�}��PG(��(w6|Y�q�$�9����Y}!�'�td��-=��	�B�3�O'W�\#+�q�O��n=���R�Q�u��{Ň��;1�^ƹ%x�t�\,�w �H�i-�bFEI��s���pfD"Pk�I��7��7��-%E�Pd���&o���t+ѹ��W�}�.��'X�_`�H��)^&S�BV�*�)[�eZ4�k���Ñ��3 ��}c�K\'�2�Rqi���R��F�)�@Ig
F-+'�HA���#k�Ⱥ�-�zaT5�j���.9�U0@X^��_-�@-��,4����~���젺�r�|e��N��p� ��m��F�H�'��oH�;1�I����`��U:�{a9\��{�;�!L�9LOv��+vWx�&/TB�3)�+��) O��M����\�?mU����h��R�����#���}0����2$��������s���������~��O>�J��8�2'�k?^{�@C�V�>$�>���i�����*\6R�#�X��5Sf�=Q U^�t6=� \�K�4UQ� ��R���@��ك�]���䡵�w�`ߠ�M��}�4��P��(��`�w#�}��pr;&�ax�;O=T�� l��ް@��C�h|&P!�X��|�p)�%@�VE��Cb�sS��$(3_.r�H+������[�,�3;�X�[&:�T0q2�L�q�s������T�`�ď�p]{�Ѯ��o�6�Ɋf��a���	����*/6�#�K�g��~�u�\g�>�U4C��L]����4b������u��b��J�.� ��B���pܢ��$0��D�&�^�^S )��d���J:��|���cͶ:k�@���E��g��[V�w���
��/��z���zS�!Z�O����
��8�(���K�0����Y�6m�04-Go�[��̸�k�`L�0���r~���?���xe�$��B���M���.-�\* ȤO�.���*I��y\����ty�r�RO�N�<}��׵���*����v�3�]Z���QT�M��5���-�cLБ�{�\ ��i*�OM����ϰ!�7�l�"��r�U�-{����Q�1ӟ� ��c�uOV�֕{j#�dP�[@�%���U��[^��u����+�%e�[#S����۷�j
����o>!γ[ao�I$�?pi��a١_2ݚF���N}A2[/�֛�	
��S6�j&�o1�(@	<@I����>���Z�A9C��G�z�6S�"(4�r�6g9��ʺ�����F&'�+�U8 ��u�^�v��hj�R'Xd[���k7<�C�y�)��]�d��u.�DAa�w�$�R(w+=,���x����6�0��]�r���Z'���� Q�!��}��ī��	2,�E�h�kX�&�=��}�����0�EP��W����P���nM�U��(�cF��]�N��w�{��鼶#,p������;�C
��Ԩm���h��~�|P�vQe���Pl��b#	70��J��_�I�����p�'
�������q��I�M��q8W�	q��rX��TZ>�kD���e,s�|>C��r�-L����T9��f��a��� ~��K4����{���}������9�������&�}��<�9�$���?���@��to*^�-7-�%{�U|D����oa���Z8G����D�A[O,|sug&�9�L�G�Х�^�����(,E#GO����¾Ԩ�t��Hᐌ�91��Opr wS���\�o���S#.�=a"+�\��n"/��n+��Ԅ��hX�F�S@g�o�u�(d�0Ԇ�2��CW�1E�<�L<�k
�BB�T����vG�F��m�E=�W�MQ�N�0�Y3��������ԫ�V��0Hѭ�;���a�D%c�g���F�-9ՠ5�]�t�b�T&�����Tcj�Ę�Ib ��u
�-��Ȑ�hD�0��|h�)Wv�Ag��-��S"A�tJ�A�#�J�\"�501�z��!�TF��m���%DY#)(�x�q�{�u�����o��/c4��@���k���)�9�T^/���h֥i�f��mѶ��Ru*���k#�(�J'r2cl���~s�I[�P^����+�)p$
��1�Р;�V���ߵT�j��z�Ȭ� �87�6�z$��ȴ�s��q9�:����uH�
jO�������{�9K�+�;��X�p�	���g�U��.ST�_�%ZZ���UH�n���cW�e󾫗8m��Hf��\��[�
��3�AxO��	��v�5�]	�1�
nWΤ�9j�m�/D�܁��cSJ(��r=4\k��0��WB|9u�Nف�!�ɖ����%ZO/�g<�69n��&�k5�R�;H[��3�MW'c�� Їl�4Q.��wv<I\���D�2�P:�������K_ˈ�j��)���yg��9���������Ǧ�^��H=�.�%�B�O�;s ?Sb���R�a>�@RQ:~�i�	�{
:T9u�&��v]��poH��a�qg�G�/q)�KBPM�[�z�j�(TOI��ƔZ(2�	��`an��<�:ʒѢ
{e�eX^�~2�O��A���?2.�7[q�#����n��
,Q�N��%$lK/	& h��`l��]�?К�߯M�E�$�R�K�C��ti%{3�U�?����t�(��H��U�f�N�Zc���1�|��;�JV�cn}�[z�s7H2ޡ�-'�ý�[OX��#�i��z��El��d���.�ax�(�W�AʋG-������e�(��1��y��\]�U��V�`�i݈�����ʀ��)��- ��;QK�K�+ؿt>�O��xDF��H�u�y�S���O���0� ����5f夿��Y����J(��L�4{��1�I�|t�^�U�F�+'j*9�e����F>��<G�Q��9#0��x1�8��21��m�<ߜW�/��)�]N!��`��! �|g�~���3Z)מ�8�X��|�^rm�[G��@Vq�
�&�7���-sB��ʄ�'K�������(Z �&-D���/��`�^*�w�?g#�d��U8r�[8ח��Bئ��#ч~9�3�Hw� Y8����!�ϴ%0Zݦ�oX��i�*��x�jk���J} hO�
03��599��vC�������܇PsO���I�H�$I�-�@��ș��cL�4�\�q���g3[BB.|)��$��(�h5+f6�H�&�~�$Ĺw90�1,j��_�VfƊ����8��Ϊ�U��@UNJ=��ty�S<�g=O�D���9��v��$O��E.cy��5��#�TF[s � �G>N��b���y!����u��5�g���ۛ�W_���U�b�o�8W��]+ �"���?&��~�?M���N�)��WI�����'g/���Ἧc(����L�8۾͏�T��e���?U�5�*�!B�qv�#	Y��N���?!'�t���Cp��9�cĘxb�e�2��}SVa��4>Q��1GΈ������E�O�ǋ����Iu8�����i���\"XF坷X��[)�&<z�'�~���yӆ��M��ɭ�k�n��\�o>kTr�HLU����\5ٰ�^͸x�3�Q6��^-r+�Z�F!�e���&�]$;�n|�P�]b
�o1J�;"��ʓ>�2��̓�z����(�v��S�ʤ=��;�Z�p��H{����Jiz�(vi�����Q<�5m�`6���MN9�g��s30�M��t�D�|t��>��(r���Ȥ��MZ|��w���J�e�>�_���
�D
?&$�>c����j	rk�~�"�quᾥ
C}@ꈧ��eEv�ۻ7/q-�)'���|pkvȹG憋D�#����������S�ނ��I������A���҄�-n�*a�%fd�\��hf�+Y�w�p �d�I�Og�����4�=v5�r�{nuX�+�y`��g��r>���HT>e{�\���h�d�ּ�i�Q���=��aM���m!�9�g�"��N��;�8�x�/�l�&E:h��UL���KQ����i�*�j���&�HЇc߽<ST+�f�Vq8B8�F=q�32G�ҩK��(>��"�{��t8�z�h�y�j�^R������Iblh������J����� nsq�e��Y_��(�R���-q��Лʅ]Qz�x����M���8X���yC���� ����%9Cο�!j�vi�aC1��-�%����2Lp!\L �Ng����~:������@D� �����NI���ѬƩ�D0�GA���z����C�痭Ω������bƶm���M�X����q�f�k��������O�n���#8V�&J��K`X<՜�u�F�~u1@
v�G��Yӽe����=_U�p�����w�M�wׅ�����ڡ�?;����oӄ��@�q�L���\2�(�Vɠxh�N|ւ��|�8��q��Jv�g�� �����G�4������3"��4�5v��L�t��f}(�y=�3z�w�	=����U��P6�,TK�}l�->�]u�y;��x�0�A�!H��Q�W�s0*��g����B�-��+�{-��>� T؜�S��/�z��!�������_�'v�
2�:Y�7k����;we�i"��l��M#�O�?���#Q/5��|!_S�J-y6-KU'���q�Y��f�?�����Tl�w����{
Ի�sTW�%V&����� ���C�$K:��V��@@�J����ϖ�e�B�n��P�0�a��$� �:�������"�f}7��҂�1[��t�34Tz�co3�k�	w�#wAd�������f<��m6��|g��j��-]�A���[���G�����4{�Y�ұu�g/8b�0ɵ�Y���˲Z��=���Z�ȹ:G�X�����~'��6������N���K]��Sڡ��)G�[�.����Tt��9�6ӸN7�P�E)8�Qk�]��^���-�H&�)>�`����O������p4�V�j\M�O��d�����N�T�|�bA�T����7̘��LDjj�1@���=�=);l�Ʊ�o����ۺ��cl�t	�B!��Ko/�n����Q|�\����*�9��Y�h�.�pZ�;!!�HA�w�B;�d,g&O+��,&q^緞4�4�|�������ͭEt�e�9t.v�A�y�1_m邬$�.:5�Ϋ�)�`�jX�ӓeߏݢ���w��%��
��u�!G<Lt�.���J��	��s �.�C�8#a	49�un<��!a�[&��e.;��k)cZGy�'h=vKe<ӳ`��T��p_i�4�|\La�G$CY��!Fm�ycѵ�"�[ڋ�{��;�p���m�7�����RX�
���p=]bA] �*^)%lm�xA��}�'5�d�#�XZ2.�9�?�K����?���U�*���J�1K{[�~�u��� -`�O���X!���XB[�mEl�4L+�)��:�~%�fs~��8����p�/ހ+��q .$�ުt��FN�Qc�e/��*�"B���Ņ	�g�U�}1qTk��Sr�N��хsA� �)Xȵ��0�8�h�����6����g����,}n?���8��j7F��j{v^7�u(��Fk��̧�la�����o0�����}:?�gހ\�v��Fh����~�D�}f�Ǎ?󬇻c�R���&�f���Nt���a	��m��@�YO����j�n6!^zA	���ݹE�y��&{�R���>U��VH����<�k�T��_j�&��Ǻ��M%뮿C}I�0����ĥ��A�I�z2H'�����6p+U���oQ�B���<;��Fu��b��Ҩ�+d�hΪ�w�<P�q�
fO'n�I@ʉ���/�6h~��-�ݕhRE,�0��X&�t�lAE�.��E��$��4/#�Q�?����/������~L��3m����?�7��+��b����2�L�0���#,�h��>W��9�荨�\����B�=��#�r��!gi������|�C�q�9�pA�F����_,�Eǆ� ���#c���7�m�̍�\�t.š_��-k{�ɓz�^g=r�Nŝ���v�||��ep̍gQA6}���۬y��]�Խ��ML��emp�
�D0�bv���Ӄ}c5C��,ՑG��+�fqs��Uof@����^��م�S+�QB:�����h����Sj��7`�0�5�[�qB�b�|�u�̖yex�������	 5����^="����S'����<K#+g����ܐ��|Bk����ʅ�!4�F��F����W��J@t �Vh�] �W�{iP�*9��!��F*�Oӽ�����?v	��{s����,w��h*���H,\��xbm���������D@S��G(�C	%�Ŧp9�O����sy�+��p����+�1�����G�!`j�;+���$z�*����!���^Q5Tk9h�-b��}*����:&�U8d� ��P���N�8�`_��S��3�H+9,��)J
�3xCW��!�ٹ��6o��>�$8Z�B�߿��~�z�������8�c_�Ǉ�B�.��A�r�Yf����)�ZǸ!�jh�\@���2Ȇu򇓱����d�=��K�2Ǵ8�ln�TҢIP\���s�����MR��h���� 1QX���	S�BW���|V ��9C���}2̥�MN�E��۫���r�ظ����Z�[����"]Ϧ{�]�6.	�w�!�xN�H��L�*��7�*�IGlx-��[iE3�S͂\�ZQt$0�S���sw6T�mqV�Ϳ��}@$�ψ���a��".K=�R�U�!1��?C����
��r>�q�3�b��-�(N�q��0U��b������qk(h�p�Є�jtU�F`�h�za5H\5�$����3���t�,|$�̹��"� �P��Av"�)��*���%?�y�����ͯ2i����|�G}Y�m��9���U%ӧ�`e��G��aZ��mG[W�n0Qq���t��v5�3��e��+��y��_�"�,kV�A,&�Â�e���kZz;���A��*�{�g�ф�.�٢��w�~\��I�i��j�Ϙ<:�\qfF�/uq�\�nՈ)�h��z��X�˕�K5����~�*�ED�r.\|v���9����돈�E�I���~ă[��W�V������X3o��#[�� :�5-�g�GL���1��#yS��Pc�t��l���f6o�,*�t[;���_��E�����V{(��?�(�Zv���� JQ'���Q������3ٳ�x��U�al<�!�<�"q�F�̙41z~f?4��
Yh$����^Z�F;K'l!NAM}z����u��:�a����q<�d��;�"���R���\���м�zyrpkڶ��B�8%Oa��[�����ʟ�Ѡ�Z@u)4��&HQ���x�z*�V���;[��35l^X�>0i�ʭ��X�T��.�kpɽ����uN��1	VSƊ�܎�=�6�G4ڰA�Gc�Y�1s�k>Aw�h�mm5Z�v��c^�:e�"�2�F6PF5�:��� �b.��AC3���```��C6���a�` �!�vw)J�:�Ô�>�!#�ɭ6���H�<�s��_�եSJ^B.&��/�ʥ눝7gO�
8�����C����?_�8�� �e@x�����8��4����1P�ߕ ͍ĩ�6����Y�]��t�]�x��s:���w�@)�;��Y��.�����yw�H��T� ��3�y��8�,Dl^��$VCV���$���d���H-@e���4$�FH/��"=���4�5�	K��:������=��Yn��3���Xw�pC���H��,)Tf�6-�K���_�B�#�6;��o���V/���_�GQ"���!=@���Y�Ū�K���t�B�ŵK�\�o|�3�A��IVˮ�D%�6*݅��$�9�Z�c4[�^�;�t4�&]7�T�pp���u�K?&*��9I+�����mgy�ΫZ1ۀ��d)���`��y�LJ"=�Z=%�c6�C�*c�@ޭ|�r�pV�`X����ݓnd0�0�V<����	����X�9��X]�^>)a�U�H(���p=L4y�B<�<ť��/(Wlm�z��z̋Ҏ�x
�f%D|ok'�y��l�������i^�À�ŗ�/�|uIRX�V�N������/�4�*��<���K!XM� 68��"�If|p�J������p��a�lt��9։Q,Θ�����U��WM�fa��$�{tK��m���/�U�,��Y�}��ZZ�q��'[m*����H��!	2��F����K{c�J�%�&ϖQ����U(�tQ��ܖ�Z�#��t^�8��1�@c��<�^�(a�Ѧ�jd���G�]�A9��3b�C#}vϢ�eD֎��~]T�&�����!��w��߮��n����%����DoK�,�s�D�g�
aU#H��Dm�Hq�_����}*�����<>�o�8jUM!�E�0 �!�E��*\Y=FQ��û�� �Po��O��؞�]v��mx�&q���@�lG�Ck<��
��ͧ8�_]}F��D�4��@d�(^�b��Є�`��AO�>�S��+~'D�6Q���1�!���*+4�Ɂ���S�}��F����đ=�C�L��91e������R	VK�D]`ի�g:�X�jO�u,���Ͳ�Q�"�E�C�4s���߶�3$5�+<��l^�A��$�����I����s�6��Dr�L�\@R	S+56�2��޹��b[��`��x��`ff����D�<r�k��V�Tܬ�
d3�/(H��fb��4�)� �kG��$Y��ˀ�(:� E(�O�tO� �@rXK
�m�*-e��ryt'pA�3%�+Y����Fǣ`�pl��f�,n(l���tgķ�*;	��k�6���^��	3�l�E�pRv�5�<�̫��i�(�-݄�[$>>�ތ2�N%��'FC�IpR��V0}��
4Yy��DȔA_ڒ�p��|�������y4R�/F�ň~�+�$<4�h�@�Ք
���Mʻ���}ѷ�Z�8�qFV��T���I��O̩�Q��+_܅�}^���d�@mĜFg��������=L��$�$���$O9���oR���q&��J,�=�9���f� -���롋�dz_���9���h0�`$��MC7����^_�Kcg+;1�D&�4����մ�anP���~.�C�ՙ�9F������nץǶ�j{���������c7���i�)J��=���K���L�N�-1ZX�P�?{^��F�!�Iз'��pY�(��ﷷ\��w�1}�	�<`�˫��d] �`ڗu�2��w�9b.}�.࿀��
�����r���%�߄z���&�7	ܳ�Ȑ����1/
�Q��%�7�GAt<�%\���SY�f��ҰJ̗m^<1�[���D������O�u�og�������;�찭�H!a�8	�Bj�S����3?c�P�y��ǉ��y�4�?6�|�x�{b@��d/0�m��z	
p�H��Vt?�%Py�e��8lTJui���m��U������MS��6� ���ivEI0<sYp�Y|C$��5���@�}�~Ň
�w�.��"!��a�w(�ؤƥ�-�H1mC</������B=M�N�a���I��i��=fRñtI��l6����_DS�0a
�&�Y��@'/J����kq��OWm;&x�;���K2�D)��8�'Sr��v�Da��5��-�R�)X� �Tώ�3Q�U�XR�e	����%]qO�����6F4�TB��t�=��eǽM��g�U���\��m[��w�V��cg 3��s-�\��G@�[(���`����+e�(2LCX�W* ��P�o�c�׬�']�2�?d���6kmV�x+D���CΏ���;�P���_ҕ�V:4H�-1ȅf��h�$�ɁD>�&�4#��۷^���`?U-��g��-؞�8u\�`�h�@��aCxs�Խ�|�j�}*��^>F"���	�������;��]�EZ/n#��;�K��Z�� �!"A���
������3K�
���z��'�,J9+���[d��^>�&��I`Mxf��b��SƘY8��s�KG�g���^��:��k6��F�"�q _�F�h3P�ʘP Č����k���U�Ԁ�c�
 ���t�,��a�T�^9�E��u6�Q�+�#q9��B�C��Nȓ��5��tBk�m��a(��T
c� �da�1PV檜��|]�nW[�!�C�Uiw��L�E�j(�e0&#��y@`�	�.-�lcq{?�1���N�Q�K�ρ`9��>�3kP���V����d�ua Us�%~lp5��i�<K~�.I(PS������+>4<��l �Ct}&(����U��i�$�9:#����-i��ȏ��8D�GD]�1�#�2�qS�AC>��0��.P��$�<Jw�Ɠ�Xcf����1�텠x��?o}����)�����}6Sz�g'�<�*̹�<%���p :]m�:�:�
_�B���30����M�9�y8 �Q;���-�"C+|?���\�Z�������<�%���,�t1��\��޵D�� �!���ҺN\��T��ǖB�����F)�, IP!R�_��Q�5�H��l��h9-eP�N�8��|������Tw �J:*�ߜ]h����z�WG��(Mr����l�|W���M�\E>a��Q�rxu�ʄZL_�y8!�6z{]��x����.}�F"}mo	�m�
���=�W,��5�ؘե���'�#x,�K�HZʟ��(��������V����@(ݤ5��h�5}��\���X���A�����ɮ�ǡ�H7��kߟ�C��U��;@S|雬1��+|������U���M� �v���g�!�����#F[t��Lv3Lʶ�m��g��!6z!�,����t|~�6>Ô8�b�����t�	DY���n��z�O��V^A��3�E %�e;1Ɋt�C}T�k�?�=k0�
��mP�ۍ��c&?E���(�-�F�J$|���o�|ȫx�!_�gv�����j�	�K)֯c��ə�Ś�բ�ң�X�'�c���	�T��ޝ�:�͡��4j����ya-:4���d� !�+���2�l�'&��o5�n�>���i~�ԁ~�	�����YW� �.n5�O}�����<@�ihdpb�����N��+#p���;����{	�4�Yu�u(|V�_XY^#�j��D5��l헵�P2A���\���G-�j��Ws����� J->e�UB���E��Z����[�����%���.L��m�����l�;v�7n�e�$�@�0�i�:�7;��8H�C�R��f@����dվΐp(�=ykGi������?�<�v�TYТ^��>�=����5��1����x�I�Ր�H�W62�2Ny��S}���ɾ��k��m�9�tdPZ���}����y���"�F�#��J8�E�7��v��5�%ŵΙx��/�ʝ[��0>��=U����%��5�M�}-)LNٰ�0���w��!�u��q4��ԕQ ���㏤Hs�v��uޢ9ˉ9�ǋ�QeZ��"���I�SY��.b{���@�'8sþ�� }Ro�F��C�T�R4�����6��"�#��j=��,!�sKz��0fP�������Dܔ��貯����fD�&;T/M?5���~�d�|��$�k.���CX1��bMt��m`�/��3e4��T�k�4M����Q^���eŘ��AOT	�=�n�faҕ� ]%��c.��AJw�V��f��|��Bmj%�Ǘ�3��ػ���'.@m�7�?��2j�;���c�\��	���Ã�Z2��s���>&���U�0I���ʿs�0\���W�I�A�0 d�ë&�r�N=_����V`�Z0��҉��\f�2j�hg%�A���J���%Ϲ�",?5�5�O���t���qJd%��M��ti�,���L�
�qPnM�#��궚��G�-D���)\�CFg��2/�=.�����n�Lp~쿭��R�ؖ�l|%�|�K�?ʪx�z�Z�[� �A�7Z��J��)q�#�Xw}�J� ��0M�,�e��{�����5�����ͷ���%l�� �M8�����|A�U��~N��`�ϟs-vjС�k7!P>S�׋�6��p��E�jW��N$tYM������v��)�U�[�ݷY���J��AB�x���Yy�9�"���҉j�΅FFn�"n}8w~<�[����10�Y���T��|gr�c/iI�󭄮2\��/e�W�˃��=�U����"�e�4F ������yG���$�`o{,_�y<��L��+!]���E��~�����Xk��CҊ�WB	@��զH�:�%r�.�Tá#�D^d���"[φ�����/ג��aH��[�L%���#}�u#<ǋ ��9��	=nHDe���B�����r\K�&A2&}��|y�d.�8ë��	d,������R��ϸAH+�8J�.p��	��Ay�x������@�D�iʹF��>|P���鋐E���r�7Ш���UVO�Lo��	LP6*	�
�7t�" T%���A@�߈�����(���>��>R�W˲�:����"x�Z�r��$&H���^�h��7,�(�`��ϋ��`����А�!�p�j<¥�szڬ	�<��V�+�8�q���G��AP�G�:P�I�Ӹ�噳�� �jD�
��0�'�ϭio�|7Ry���Bo��-r�'���Oǡ�<lM�\^���zx׃��UW��5���s
J:!D߃�����~���|q')y�g\ۙ���8|$�r�Z�4)}��yI�������c�f��v&YB��_�SN]Sj/���F��#�[�).SqƏ�\����l�����/��]���]i�`f�(E��N���+Ӗ�{��f��47�L��τ~~H���<�<���4a�(��9�5����2�����}��G��Hй��l�4�oH������u1#�N�b�ld�N��=WU���-;����8��W��*u���L�5�.�;�9E<�q�A¿�=s(�mA;���.����3]��U��R�x4ך.�Y�),,�"������C�نЏH�\���n���@��o�<!�$��jBM��(a�/�Zi$����iJ�6y{G�y8XvHa���}X�:�smׂqH����-��;��|!(5���R�a�
-7��Q������Ky9�4��%��k_��X�9>�
�&�l��J��{rtQqa�"2:p�m>ˍOXu�
-�V�\�I`!��umH���J�b�#c8]�d�UmԱ�d�[��#=��kgi���2�1燏�D8�B+3�����y��TO6�]�u�ڧ��=*�Zc��^���C;����9%�b�����@��	[]	p��y���z���H琸�N�w�QRg����f�(É��<�Ǩd̪r��t�A�\?U\Ϗ�1`i�D0 &PSh��γ!&�mft�1�6m�O&���@��������^���4pl���!bU�VE��p�*���d��56� ���&����2���y�Gd�}/ť����~#��I��)��>k%r�bD��
�t�~����ľ��T��J1�v�Гw{TNQ�w]�4�+������TvQj�n,�c��"?�'4.����2cA�9��\��vݙ��a���z!ȂsL��_���G��.�BՄ��DxHF�	F����p�df�o�u�a��$
/ssg�0b�E�
�@�Y��|��Z�d����C8,��
5�˷sS�|�Q���Q6)�!��N,��,5PlMp�A�A�Ħd��j@�)-V#�'3��;�$:��{�_��i�ټ`O/���F�T�Q��ya��IZ�`!-ZxO�d~Yɛh��c��=�z�G�"���~]}۩Xp��k��9�J#�i��N!5�aG�ʎB���]��Dr�#����g�i
��7�a�j�@��!ʑ��䚠�͌v�� GU,���Bj�V�&Ei"�`�+f|[bb�`����.�@��)�,hȲ�ʽ1�
L�8am:�Zl���b5��b������ŵt��F4B��p��U��\"+b�E:����[���ߖ%#�Jz7��|>�gu��?GW�r087ek�������q*�v�\��8�}R�vsɐ�|g��	�6��$����y�{��y3����kŘ~/��1�J���r�J��h�Lk݀��W�/�md�-�h��@hTA1�p�Rl��}�R�p�
)N~ ���`���>G��7���٫S�H�eS�e;��� zL��e6��\���A��Ji�E�B�I�P S:�5uaufIlUp�n^٫ЈG���D��x(����~�x�9I�~;NI���Ms� �7���o)�'�$ƍ9J�/�Ae�-������tv��b>S  7B�~et�p��꒼9�l�|�R���J��O���x��M�
.��[qWz�v_,ju5D��ew.��K~�o�X >�
��i?�#��y��󡧡��e�;�p���Mm�M[�^l.47���J�8���U�H�k��(����dSC�0E9a�
C�
�~���\�ǲA-�o<� ��k�lrM����U��R� �p	-!�Q���0Τ�M�9i�­�	ϐ���0h+�|&�G}��d�B�8.��� �U6��w��$Dj:�=�兰��{�?�K�yHK�Is%��nJFΌ���b|�ݳɐ���BI�uo��T���Z\�cB��Kg�[aU�*j�jkZ�6 b����&�d҇����FEۦ�5��ln��d6�fO�%K+�er�V!�/����4/k_��?�Oj����1\����͜w��K�x.��K{����2���X7��@O>�u�,���e����-�ZZRi�~�Ꮸ�0�^Sz';r���������M<I���Q"~��B-���"]�K�-�J�],��nn=���GO��n!��輓B`T��e��#��z��[=����ef~j��r�#ǳ|0�������t���`jnE�3��H��a�@<U-א�nQ�?�`�n�3OҀ��)���M�*'�Uw���<��v��%���߰l=��V��#�*|�ۑR?i,J���l�)��G��/\����`����T�Eg���{N\]X]�M��(0��a?8m�|ݍy\��a�0�5V�$-���t|�׾�v��E�'���G�D����T�E�aLCA���%�=������,�@�V��h��lU��z�H�!!��,��-�_����*�$��U� ����h��Mi�"R�x�uT�#�O�ݞ:�K��r9r��BR�7\�I)��u{��g�τÿ!�Y�Ћ�$�-@ށX\E��>D�_0���v�Rs�V)��B��CK���µ��D�]��=��gTY�J�7�@�u��'(:R����%^n��"Kv�cr#�K����12�L�t &�i�̫�΢���s蠦aV-�K��Rxʲ��֊�JԘ,����;�:6��Њ�G�m4�K��?|�D4�3~=�B�����[�X>�e�|Lu֤@�VEd(��\у�� W
8wo��^�����k����z@8wۧ�R$��kʴ��@_���]�EB��2ƻRV���'�db
���[����歝m�8���OQ����=Z[(a�4>����+��{�G����I/2����/�)҉}.e����#��+���U�_��e��%��[p�2ik���=��7���Y�u����<�_⠊�����0�Y*�L٨4�+���N{�5[Iz+9���x G0�YQ J�ָ1��CG�mYa��7�d��o�V]�tz�l�#^l�S��M�?&FJ���E~7/*��דVn�z��űO��_�����6�4��-y�{\���p��1^��a��#�Tm_Ikw<nA6�Or\��8GYr�*�k�q�����f*�~^`E ���m����JS�;��*W�1XMb���r�6��:G�C��U۱�lԔ�0��(ɝmP�F��;�fQ���,��tB�ܩ8mm�^LR�}��A>�c�A	���?M�?�[�:�HB������Qҝ��ޠd�Ti�1?��-n�-�f���������k���%���j�� Zo�ۚ�~B�jMz��E���8�����Lܗ�c���4�ʆeV��dn�.�)�^�~�3kz-Ru|����:�T9ȝ͋F.�Q�B�`�0�S?M+/*x~u��T�DS*Z�v]��t�m�jl 04��ރJ8Q5�ih�3�+�(�ҺE���L��W����Խ�a��D���)�U��2b�v�����|xFM��w��bD6l��J
*3xh^7��j�7�����X�� �] \��ۚ�]g��tUb*YӨ�|�{�WJa�����vY�b�� "��'8��KZ����^���=�8��#U_��D�E6�g�<ì�4�����4��54y��<�������zh�˒�r]Fx���+i��%�	2��5�k���8LfZ���p���y�n�<0���o�P{����z����g�X���.�pS��?�w��wS�+�ւ9h��́G�V8�p�eAf�QN�p��ƺ��ukc�g~�!�����6I��H�����#��"��� ��ᘲ�L��1d��q7���k����>끷���
�A�CIG.�g0G3��g�?���m�m�o��i��QK����Qb�&e���VS]޶���iWE��"F��?EW����2�R�!���A�U�S���c6��f�s�&+����}4!�z�*��y	K(T�Ł��n��DTD�^�%����$@�1E��wM]��k
5;�>�+?��f��9p5�K��	��� �Zq�f��ٿY}Oq������]��ILʖ���4��I?^�"C���t��\�o;�8���Cs�ǳA�<w�j|��N�b��k�U�:(X��m:��:X��VK[@�����}7���W��Ϭ)��I냸|E@�O6:��.@*N�s�0ż�Z�����x,�䆼��
/���鰮�1��E�d��\����!�i1��|u�p��;z{s�ܧ鋓x���n����SϹjȝ�] 72�F� ��{�n�ܷۘ�&�L��@G<�o;��H���`7��p�sӤZPx`%� 5�8v���4|3SW���}�t�̦�N���}g�Ba�V�R�P�gl�u�2ٹ?6(���g.�?|���ML-��&�!}���]�����&Q�֘�6-6h�Qq�o#��(OUҰgҾ�P"KQ�ng*����jU���[�1�rj~��-�4◄�ya�;4��k�#$Dۜv����q��L(�9i~`�P�yJVZ�R[���!�~b�=�Ʌ��$�ۻ�O��A�6��j2,i�m���M����]]c#$��#���Ψ|*����[E�������-�A�1vS��ν��k#�p���a�&U��aX��ݠAK��h��6�3�
ޫ�p��r~4p�/�)�h}h�&�|L�]Ƥ=�ft��[M�����t%���v[��l�mqb���:H��NX���1���E�w�S� ��Uwm(��)Ǐ�bhe���M�<o�^;'{���A���^J��;o�z}�0Q�g���8UU�����{�o�lNA�Gr����6��w,�˒�ɸ���~B�Ұ�m��-|���6�~j���g�Q@ӞQt�h77�4�kf�
O���6�����J[
�$�YK�R���������c�����3Œ�m�4������ߩ[(2V)�X|}�#�	��BŨt����B�=_�tҵD,��Z�ʪ��x����lQ�z��&hS�ì��w�^A��/[BD�K��V�1�,�+=�ES"s����׻�)��5ҩ���bAK_�FƧɊ�"C��[\��]R�Q�>�������%�w�"�ߚ�����7xe9!�����p�Kvf%�I�pb R�0f��t�ĩ��S}����\�^jS������:�D�\���&��?p��wA��n��gII��܊��-��H� Y�r�'d�*i�(kew֕�&��s�g��l]�&#3M��c)�*ػ��|�"@'J�(���!����V\����f��`~�G��ů�!��Ix^�˹�
����2���L[�)�w�c���#�L��$$,Q�y<��-"�D�#]�_g�dV+�I+,�G��]L��^���W
R��~���9��`n�]!I�4A��;홎7&�Pke��L��g�,hM̭G�
f/��J�#���NK�?�ZO�~�QΏ�����4h&�*L_dv�Q�"��zq:Wq:�4�Ny�� CW1�Nw�Hcq�� ���a@���Di]X���ޛ�>9ïa򎼾��6��V
�A(`ǉ<��%��Y���۟�G��.��q.0;�&��~f�osm��Y�|3�|�]	OX����	������H�xC��p',�r�t :����`[h(~��^B�ck��~̡\/��荼3����-ˌ����/l�Sn���ڬ��
:��-�Y�dGP��>�o���<!������o�gU:V�4a��3��AJ�����f�)nm��Q�Qi��2�օ������z�$�}�����$:}����ܾ�/������v�s����Ď3��[G��Y�q�u�����,��q"T6��Cj:��fOC��zn�	ĸ*�{�x��ѯ��xJ�������U�<�}��5 ��=�W�^���m�_wdb�L|��h���O"`kHSA|z/`�`��I�Xs�!#�P�o���.�ܫr��xI���$��"��5F|q����i�S=�N��&;Q�-�b8���(վR�R8���Q����v�-�����[����R�f�L1�.y�Kē�r1�IM`,������r���7��L�b,Ġ�yu�|ǫ	���{�|��qM{��-���Ǧ���I+��U���bMq�e�xϢ!6�g�)�� ���>�9��n�]��R��n.� ��u���ze�n.����J����u���']��ޜ��ȫb�8)#XL�x��_����(� �V��pU�]������3�R�FL_��mDQ�w��	[�d�7�����!�p
P����g�|Zv�%�A:u��O��0�b���)#����U�˛�YQi[-�$�u��=�G|��r�OSbK��^�����Dq���S�5W�l�m4/��ۖ��� ���_=:����`�z��kEOTͣ�ӌ͒F�h�p��	W�PjD�����0oݯ~ۗ��>ZX�:�Ί��&�*&�_��X���Z��V:{�tXӰU�Ș���P[$J"���lN�R�<�U�L=5'(� �>�a�i�Kew�H�.�Q^c����D���O������%ȗ���Aq�^�ξb�!�Nb����*͙�k�:hL���l|c}V*0+I;q���T%�݂�vm���% �r��g����[4	�4���Ķ�4we(�g��Ƚҥ��X�'=�|���W����ĻG���ͼי�p�ф�
~���a�8k��gG�Ez��h�V��}�K|{���t����6�_O$�cn��(��o
����i�6���jI��vi�D3Q�0�iT �8�A܏��� y3���*�ϟl>m��|��|)�~�L�V��6��k���s<�qp�X��e~�BW|a��j��N��N��JK\%� �Gq���JKAL�;�����%?����:��*�A��_F+�w�\�e%�f�	4�)EG3k�g��u�3�\7�Z��o���`�=@�ߞ�Ҝ_�h��}�������
��j;v�T9�� h\N���ͦ��b�&� ������J�@6��Y�[b�x�e��`w�8.�g�+��N�ޡi�����S�$��OЌpM��5�i�y�9�ET.WW�gr�鎛 �������dA�R�冼�vh&ȓ�#)��"}w�O|�^>���N�og��������dl����������� ��؝C�`�-*n��Nξ��ۅ���kf���S
B�Dzly��bq�.Y�vNQ��?���d�c7��Y�^�ݹ��S}��M�o<��� P �ԒSVl�"!T%�̖�/��0�mO\bӭ�}"	r�y�
�{��Шe~��DY�'Lm�d�,�f���?���z��T�%��Rg���e���U�� �S�Ss�X����S�Ҭ�8hr�B��1C<1]�����I�q4 B����r$��*�!��g�S���4���X,ρB֎���܏�,���~Qr��g^ۮ_���1h�[���q����R6�6��i:I���_7����������ni�Rr��Z��Q������V%�v��+W��m��V��bT v��c�O���y�=���75ZA�@-�qoh��w�?��Aû�k��ǐ�X�\=�
8����fWU�I��AR�p���V7Ѷv/�Q�斩���Ȟ���X7g�ݡ���(��ez��j������5���'v�C1�Y'�;;ۈ�[n�|>D6�UNeY�Q��1W�FJ\.���C�r7|���>/��vח�+�(5�D;�9E�1�~��X��ݟ�&����]Ic��aP�"�P�@�4��
�&�^9����O���N�p�|D�x�k��f�O*J�qm̟*�	c���c����
���ɝo�}8�v���n�s�'R�6�Xp�d����3=XA,W��k��L��c�R����lZc�e�s�f(m�.�a���a��*��_��5��D�kpw�8I��(�SZ��	�� �cW�h��w�,f���x��`�Zt:v��3����=w?*�a�f ������ �;��\�=�}H��ң��hg�	�I5�9[��%Q�.qu'�{��U�1�3�ڝ��F�u�[��z��j�T�4�j�v/H'$�r����j7����8��YJ(��
L_	�3%�'�����c�?
ڌ}U�	�"7��@)e���A���ФA����0	�҂�y_�Hl�E���p�п�X2n\6�A��3$ >�	;���*���`Y�f�_��WvY��"m&��\Z ��w����1��`�Ip�A�!�#�>mܺ��Zr�NwG7Fy�'��?�4�GZY���:�X�C���'Isųm���HR��s��x����K����t\�!�
�i#�:���d��v��G'֪�����[�ć@�瑋�J�cwCCq8�1����@���	{SNв��^K�{��-ǘ��J���雳X�,C~���q�9u���t��f	4sj���K� �f[t"2=����)DRDM�"��]����5A]���z����L$�;/����~��?G�?#ĝZyS{%d���s��|+0ĳ���M�	�3t��[��I?�Q�#<�6���غU��_ٗSֈ���f0�1�V#�F��� ��������q�<r�C�5�Y;C��Q�<*��y���y��̌Ǔ�+��EK���2k5C/T�LP-�$�-��zN��*�u����g�'�>:�I�ӟ�6gQ�UC��[��rGn˔I~܈���t�&�'�C�����[.DI�����O�r��KUjVI6��͍����E�M�(Eb��&S�����|�3��pX<��9��n�'�0��E�C�g	�`;y1�Yʌ�P�b��p2�a�ےc=���u�'j�J�3�A�S(~z���(h��d'��/]I���-Op�v�%�av�Ϣ\�2l����i������vh�ɭl��q<�~R�G�(�RB��,��~)����'����g�i&�oO((�uf�W��	׿�ά��>���	�H��Uר+��~���ޣ楱k��D��z�+�~S|_��U��Z�-H`���w��g�3m<A�8Ϲ<�S��XW��Z��p'kI_��/~��<��>�.b�`75�L����ė�?������4p�O�W�&���?l�ѕh.��/�ָS�oyg+��4�{�Ջ�/���m"����N�#ss�o2=�ڞʫ����]<$�}{5�g$��(
۵��th�I��h7d"ai�s�đl���f��1)�(Z/����N�r����i_R�3>�����%�]S{�n?�����G6�z��ֽ<@LK7D���m����U�!D?"�lZyi�^�2��(gY�Ht����e�3f����50��۞ېYbMO ����V2��)`���N�M�V�i���:q@�kxK)׏E����^Pf�9���ԛ�D����Ϟ98r���@�R`j�7 ��P��2�zz6;�j��y�J�ƙ��;�4�!�m�� �0q��6{F�i��'Em�g�R�|�0��֘���O���n�E⼇&~|���
B�.��Ų��Ia޴�/�zcdU�tQ�G����� ���P��:��4��Q�sN�DX#4Wbn*�Q]�j���`V<�U�]$��	��Rn�?�A�4���)ΐ��5�%�>�ͦYYj���]��5���*�H�V����ÞV��ߖ�gULmu�{��b���o,�0'<vƴ�}_?j)d�
A� 1��ʒ���
O��W��1oOb�Xi ɨS�a�'�wD�+��!2�@Ҡ3��7p F��Ǣ'�|mF��\�̢7��$�#< @g�_:��,�NX��d��R�3=^	@V@1�[lNm�z�@.����*u�C`ӑm�1��H�C��!���4XS0s�t�d�:�Y@b5�.
OIo�,U��nLL�c�F���߾&v�f� ٶ��w��4�nڸ����z��͆J�_���/��� e�;E��b=�[���@��7J��@�A�Yťn�x�J)=j��I���L(M��*6��h�L���=�٬��Q�n|�m��i��ގ=���X��]�I��/��A��C��2����t��y���r8��o�
�vJ膸z�L��y���A�DJ3}$�9Z�^2F���J$����^�ev�Q�ɦ��f�bǸX.�t�����b?nA���b;��#�v!gq�t�4{�2ս���F�ʎ.Ⱦ�T�L��]uO�4|�U��Io#�d�f��}�\�BLv!���G��S��eG-�y�1���+�>��<���?Q`�?'@�:0�4D���j��+&@ Lɿ`x�jj�K,#�0�Q�D~�n���HVWĻ�j��tD��gN2� �(41�H�X��S��K[��1�Jn J�tV��`C;�[ˌ�>wgn3��X��N3�^������0vyG)h��~F������|�[R��\Oއ��x����+@�M��y"������v�6D�@%x}i��PF��N��rDBW�=[�A(�B�	���W�+�lk:JG'�
��]�GW^r� }��D�_)o�.�[�:��d��Y�ܻe$�K�Bm4b�����R�7�>c{���"z��n�L�M�Z�zSOԟ��(p�5%<	V��*<ܵX};z��a�y V����I	i!���'n��iZ��_���V����P�ຫ4��Fj�= AE�q'V���d89�ߋ@OR�7��_�^����D|}$�D+�s�m��h�_"����}�|k,m�Lq><A�]Y����2�m֒T�(yX9@��e-�|!s]��./V�[�W~�#�jA��i�З{N�{;#F��'(�)�q֫�:�39\۴К���xv��Z����/��Z��g����+_^
ȍ����h-�B���
�������nbsٺ!�������T������Tr���)ܬ�)�F�����k�^�S��}E��«XN5Gz��@��q*�#�s��{�|���Cl� k����|r)��DzC�|��Y�-u_��6����������� ŗK,���c�T"��x��.�\L�-��5����;?�A��|�R��}�cϓM;r�����#��JR����ȧ�Xj~_r�ńKqe��9�4U���r�ct�DZ_��rם4.��ة�L�}�6	�4�I<�3g���+�m��&ɰ[���S��Zz�_Jj]��pA��$����ҋt��p�c]5󥜪pl��u��;�q�Er��n�G��Q���T�k}���
¯7��O�\�'A�B�t�d]�Y�2��<W��a86*�ȯ55�G�p��ڝn4o�L����vӰ��$Xm3���_)��"���\�Gp���%Z�H�`z�,��Y�)�-~�s�� 4,�*;hH�~!m:�p٭��gJhZ����%>),kn��Ǩ�S�����u�S��愇�w� �B�)��2������ DjF��=g��⫀�����.�3����D_L�
xf�ϊ`A�k�o_"a���y�~��<��,n-n�����..�,��\Ԗ��%���9BQ�� �?�EUʓ����f����kP�{w����p�N�ՓC������&�׻c�س������>7�-��ڐc��6��Άv���WK<6U Ш9N�5�Yڪ~��6�E�ݸ�I�/ݶ�iɑ*qm�=��dT�k��c��O|�;#7����RR�@4aE�n�g���vǤ� �*��1���J�S�כ�Ņf�1Y�
j�&F�d� :j�ܭ���|eFj~���Be� ��D2'~������¨"�Ƨ��Iذ�*�U���B>b����t�f�.Y���s��zI�H��2����i��5/�hpF5���~���K�0��ʊ�>�Զ�j��J�J�k���S�Fr��8g���-�v���&�h{��"���;�$�Uq7�#7��]��zM��Id6P.;Z���oԏI@ݒ���%�/��V�ޮ���NU��c�/����n��3�#����qw`�'sF9�ң�"_��w�	&K��PD���fUn&��
p�WJ��l�!�q�x<�cIPW>�⚮��v-<l�*��}�Zv���%ח��F,;l]�v�>�̈́���I��%:.��0�B�yx���;F�o%3fk��Q�f���,r�~TK�=��^Q�M�"�­k�ᴑ�k�+�J#�sǱ�!�����MjBw���x�<sZ���W��Gj�y� ��䐤�@�|���؋�3�Z�M���~�:#sȧ���f�ϊ��H��>��ڭB{��Y9��
A�?�?�-�/�[��hO.벉U���1A)�&V!�J�9�E�(�]�P�cT "M|ݨ_���tn���"�w-��t�vT��Ƶ���e��㳠x�4E��}���{c�ڡ����'obp�x��
LOk�ξ6��\�8�g@��JHU�f�K(0n�a��]�}�a����t����)SV,*��^�f8���&�}�ipH ��7.�z��������/\ʷ�\B1Y�nn� `_��zڏP�8�v�܍髨S�Y?�"-�5D2JUJ�����kp�[Ihd���c�*`��J�9���
zj2VL�A��P�¶�wg���	h������A�ʼ=�l��	8�����$7o "d�5w��5��mە�O?@��M��lzk��n F�?ʙ�o�:hV)�������CXz�[{@�/�I�v�6�D�4¼�i�F����m�j1�*ނn<UP sx�3�a�S�4j%��8�j�D���-�a6�4��~�#�ø;�� uzC�8������C�ٍ�0-T�tZ´�40�mqj��n��_� �zLk+|�����x<A��|>�WN�t�t`��@��Q#[�I��� eZ�>T�W']��\>�;9�P��(���m��<������%�����"l�����B*�?�]���Ƶ�DO�־�4�7�3�p�����vD��5�+I�'��F��r��Ę�N�B�b��g�~���3��"3d�T����LF�̶�WnUz�r�pb��! ���,'o`h�P+פ���8�[�qۙ��7	cZ$�'z�S�,�t��1�	�[���dWi?Q����P�T�>��R������0���E�94�$	�g��ⷢ������^���N5�H��PR�� �>�/���ؙ&�f=C��~6|��#�K�4fv�H��ͺzLD�)�k�A�P����-`$Ğ�g�(:t,�D2��5A�%�!<�T�`��YJ92/�*oJ;�$��Oё���������
E�^*�4��Z�%��zIۂ$����!f�H�ca�n���Dց�\N8��G�2gđj�]]^FT�7�r���o�)�UG��>�Q���JE���AC��F~�E�|��{�<�����h�O���2�W�"mB�%WY��l�`�e$scv%7�k��L�ܴ����D� r�S�B$�PZ��|.];�ǹ������x���GT#1��jy��!�[jd� �aI4���F�*ՏU�[+�dsU�9L������qFJ�}y���+u�w넉0l��T���r��-,鐬�/�zݝ� ��a��1��J �y��Ly	�f����ܘ�V�W�^��E2L������E�@E���G�y}弰Tާa�9sTe��{R�i�����x��%`�lѕ#�=�T$|��pDJ��3�㱆2M�N��,	�p�U.M�d7ǯPr��rb>1��������v��i�a�$^��r��W�_�3Ѕs$�:5��]��Q��U�*=����7���ʿ�2�@�e����ؿLW̴���@Ga:*�k	�r������*�?#rK-�R��2<�g�l��c�mk�tP���h;ϫ��`L�eK�G����p�e,��sg��ւ�y�c��8bz�:%�FF3 ���<�q>�����0i�C��U�(\�F�(���(���v3tK�u��C�k�`�teJ��I�T�и�
D��U[ս�C����v˨f�gg�<OI�P��F��&J�$��I����s(^��tIw�?j�h�EA�J#m8��b�@[P��r~$7��.k"�_�L�̈́��o��1yY3#'.{��f�7���ے��Ɪ�]!��7
oK2p}}�nت%�ɒ�Y���a�xd��ΰ
���=�т�*��K8���'Z��/��ɻ�m�� L�T�ߣ��٬�G�����ceH��Vv�8]�1AX���	��[�i��ߚ���.��+e���+h�����F�f��õ��gz�#�lK;�;ُ����:>n-���)3���=ö��̿�<�.g�<s�W�Q"S��GT\�����Y�sF�C*��3��m���+�B��4�u=�I�W>��}�`�����(7a�������	��BU{^��5�����|A��O$6����d@���ռ��F0Y�W�o���rj��O�9�L� ���n�� ��2P�%�RM\��z�JA��$���-��(�	��ೇ�_	�d|��&9ޑ\����9(w�~kn��;zS���n���Ɍ�0~3h +��-RB_e��$�`���e�nnp�V���[�<Ϥ���Or�8�%�t���҆�v֤o0|$���_c�5�mH8J�a�#=NF�5��`�s옯9RZ��B���s�����⍿�'����V���Aol�K'�0�C�?_�J��}��Ps�U�Ұ&.�e����`��6�("�w=���uh�a��G���QZ�����O�����D��H��ݨ*;�1���T�Q�b�<�z�[l�iC�80n����>Q^�s��+M�M$N�1)�4�d?f�w)��8��d�gi�̫;�i|4�%�䏆ƫ-M/�i�f3w�F�@uxy���鷺���h�I'��E�Lqn����\����Cl���m9�n��@E�a��B���Gnm�rl�6۽�~N�k��)P��������p6*1D�h��л���_10���v�+l�CZ1��l$-�P	1l>q���Eo$@4�B�A�ȆKZ���`-	��RS!����?�o}#� ι�x6\�k��!�\)=��~�C�q�y��o$�o�2#�X;~\JV�ȸ��$��� ��y�.�" �>���Z�QOVJ2���MQ�Ѐzv05t��w\>�X���8�5x5��nf��S�%��kA��b���^�g���Yk]����3v7����gL�W���Z@��Q�uk�4�d|C4��:�{3�aː���,��a�f*�m��c[��b�Sg��>�-�	��stH��R��pǡ�ۗ��������	��;�A�c:WCW�7D���V��}�����U�b+L��5L���jL|��@R� �e�(��'�%@�=��d�B*\�����#����wY��r|N
���-���(�������P��� 5�2e�t����,0�
�S��wM�d�:�׃�B�^�
�_�a�u0҅v�����)�j�Z(FLN��o�,�;9a��F�
^���ny,�v^���bI�G�k�!TA��+?wʎ��LG|�ȩ��\إ�{ݮ��x�=JH�:>���Jվm�Ѣ$�LCӝ���Fc���)k��Da̒���@��gW�O�Bs'�7c6��PHA#��@��#�%�S��9���vI�'s��9�S��	Z	�`�I��ʬwJg���FЅ3�r-A��DA�R�-4�-�zP6n-�Й �	�7�(�#�#xS>5C`�9��R����1�mX�j�!Rbew��3�!�*��;�;�����-��n��*�m�&צ5;^����k��L�}�XnloO�j�IM\� ��K݇������	�����x�V��ݒ	_.��	*����:�*�sͨ���Nؚ�U��,�suA_������e_oRyf���gdX�_��t�N���P(kK4.@d�'�z��<3�1�,B.�r^��B����a��b ����N+�`���ܲ!c�u��g�P�M��a��������9�Y��y� ��BX���e���ժ��z��~��c��G�5�{�j���t#Ow*���,�<���o�)��,��d�L�?��b��A���7(�9�� �Gt�#� ;�{p�:��hda�s���b�[���ƺf���P�0�rO��K��9E��x�&���N.sw�i�/<���(Ss;���2��H>%z?�򤮇AP$W�|���c7�N��K!��
���W��Q3���E*3�O+B9��ԯ8�cf�r�v^z��g��N�8�~+ep��Ug�ױ3[�����)��.a'�!4��������Bتy�}˲�;Cx�-m[�)kLF>�5����jЊv��O�������h3��c����d����Q���(	��8�$��_n�N�Kc�m��R\ߎ���>�[$��8 ����ËL����7=]��a�#�%/
ȓ�<>e�v�e���*�R����$�Dd=d�/�-�Ff�y��r�����p�gP��ǓNU:����cufʷN�#��n`WŧR9-�E},��6?����-;���^=�Zb�G�5��㦱����i���-@�T����,�wǯ���ڙ��8���	fr�����L��[��H^�����OG��I�c[<�֋T�����Q�7pݥ��܁ʶ�ug������kβ�׭'6,��)��� G�Ue�:�VP�(<Q����`��%����������,!ج�LscĠ�c���we�5�K{��V��.INQq��y2�Q��������}�I*$6�ͪ8?�й���1c00���s�Յ2d#���@9�~G�O��6����Bр�n�?'^<aͧ��0�����ŰK���I�/��R11�H�Ѱ~q=E�����ں��Nw�J���?��ć��R�%*c:BjH��Ғ�u�:�/�Fp�4g��f4x�=n�rT��b�i5<�����
/��n�\Ba]h��9�L�[ƑH��+���9�=	8"�pGG�V�b�<��3NڕZ�����ϗ[�"Of�PL������X��kW���F�޿���򢢥� �Ђ�ҵs{r~>Z!%��\Zg�f9�Y��= ��m���\��DxI�)�
ƅ��$6-H�/ɉ��TO!��A4V��CL�M�w^��3���[��%Z���
i}8��>�Aƪ��{�H�|jp��#Raݡ����|��)����֌%��=�g|��e# \�f�1��|^��̑��qlOf-�U���"���)�_�`��-@ƅ���;���=݆i��Ep��#������A�j0�7�ϰOQ��iG��_G!��,���A1�Zr����-Z왑>�8�����w�W}O��5���k���������k,^ON�-d8	Ry�b��21y��5��y"�~G��E9�ާms�x@��0����Q�Q)9#A��vkۼe�TѰ�x-;�JQu6r�%�ȍ</�ɥ����פ��_�o�ݶp�ɓ�pP�� Ø=��CM�
����WF�݅��#���ک�s��աM{/6:'K��,��i%���2w�]���78@����E�"�dʖ�n{�Z5�(2��wP|��]\��PV�@n��b��� 5�A����yCULZ˵D
nΤ�#N3����������p)G����� ŝ���K�^~q2�u�BًBZ����2�ο�m��?(u-�ERK���g�8���L���F��crO~~�o�ڄYBF0,-�}r��p:�p$[QH�std锧�IB�E���SFz�L���s���s��3~�cL<"��EJ�M%p��t,����k@���@;��C]/��iO�T0����9��,db��YFnt>~6�`}��Q��B���j�Mۢ���XǛ���֜�ԌE�K�%3��l�B�F,xT�-Vԏ��E��`Ҵ5�OG�$��;j��-�ݏ�\��.G7�����W2U^�8a3k�{���V1�y�A_R�wc����!�xq��Q�����i�?�߆���{ &���z~]�hm>�-%�_|:s�����=����6�Y�����j��*i1���뼿E�x��z�_sV���wgy��]��YL�6�n�}�22�~RDe8�:j�|�����,�`�+�� �V~�e�z��d����Tr��s����-v&�;�3�? ���!-k�A�f����f	&`�r�h�����8Z��}��#b����Z��н9t�2^v[�O�3��zZ�#��M�q`�9zO<\�@׀@"�ϰV�KIG�Dt�������R��175����i�4�j	�B�0�Z����(����Q#�D�މ�m�W"N�4��Ⱊ2.}��$�����=�7@�׹I>�kI>?.��+�I��d�t�e�ȵ��Ccs@���a���l�#�������F�A��x����;�ڋF��^^�{�³~�	K���a%��;������"^��_����/���Z��
�X��Y�巡����Ж��vC��t7�(�����p7ׁ�eW����z#������vD�z��G�2	S��dTH:��b�u�ê��0�z�n���C۩�,�����Ēj�C�ʛT��`W��"�GU��s&����(�GO�ۡ��C_�&Չc���f���Y`'�ة�����z�.r��=�rI��D��Θ&��@E@77���mjD�`7S5�W~���H<z�H9GHp��UÈ��U"��w&�dHYu���oVZD0:ۛ�s�S��ag��ۘ�XTNe&��C��E߾)��C6BH�H�U����g��a�F����7��q�ݦl��i>r�+�]��	�5�ݕ�vT"����Q@�lgd9݀�F���6N��f���y)�U����	@�وc�ۋ��ƭ���k
I2��M&�gngV�w���0Ԇ+���j��b�J^��I��y�����}�^ZH�l@�X�􎄫��-D@�Q/�94Nqlf�`n)��f���e��bQQ�9�e�t���޺J�PE�0�+!����
Vƌ}W!}m/ձ�E����b¡�/����u�`\����N𯐽{�8����pQx�uh�R��-,M�X�d�������6��S<o��	%�ܒ[�0pHP�
����.i�o��ЧtŞ��m�IO�S��+{d:H瘽f���qd�ȶ�꫙O����F�]�����[А���c�wB��lT�2;/=�c�Kn[1��%��%*���"i�W���u��,ի��%�AOK��ޝi�T�  ��< ��A��X9T�泗�*I�%�v�ǮŪ��~!��;��8.ޜ��Ԑ��AۀЅMz�ci5�(��<�Yu&�)�m�V�~��գ:K�>R�8��/�l?���]{���7w�ǋ^ jה���>�?+��>�8e���n�N$�����=-�WhD��]��ꄵ�0N�v�bo�27��z�zy-���oQ���n�	�Ҁ4�I�	ܲz۳&�|q��d�E��Ǖ�����#�c�r4bx��g��5�$La �p��0�%�����^o|��j��.���ʟ/�1�6�ˉ/���R�_�9k�e�b��΀��F��)f����J鯓�pm�=I@��w9}/��~�N�����K�C���j��R�$�ܡ��r!�鮁ν�m������BD���\DS����G��*H��?�k-~�YR��Q{��:�%��Z�>�\ލ�Ic;h��[<�:p0�T-�L�÷*�����ܲ�� xR��Љ�q����fͱ���g@`�%�a$��N�bD�$�kgT�I�Q�~�Y�Pn}dI�ލ��u�6���zuB�1�֌��`FՆ_��/x~%aJ���t�=7-�5���T�P��Ӝ����nm2�U�7ځ��&��u�%�ݦT����t�v��F�����H]��Uq�urN: |@b������yl2o/�^�>G�[�Z�%��x������V�QK��/�F�gR�M��M�SK�P)�ú����]�C/������6�3�������4:e*�ZP�ք��;��4���|,墊,���3fVV�<�N�g7�X�e��ᙾ<���)\)s����N��;\��䮀	�v��L����<�n���&��&����=P��|�)-W��o.��n��.e�O��@�N���\�J���;9������Z��Z��v���bĴ�����|pvE��MsA�.��6�=!��+��HaSI�V�,|h�Ң�f`%Yj���ȵ�'Pg�[p&�k�}�A��x^Mb-����-8�A};V_��[O��p�5��2WĮ��R1�V��0�Ơ_ۻ����,O}�v��!DX��'[OOt���'�c�#tV��O��Rh��@�7;�{��רT�P)D��uDѐ�bk?ָ���c��م��T��rJ�*��2�_f��9&P4"7�e,w�&��]�:��bLM��С���9Ӝ�9���z/e�D��,k�G��J��ʛERlx���L�q�|�����
A�-le�q"?t��oLϼNɶ�Υ��+P�p!B�\09��TZ�T�9�#SXV�F<����\��H�3^�:��ida��IQ7�|��ك����6s�p�
٩��.s�4�FـU���a�q�C�?x�"r=���P�`/.]���Tg��Դ+݁�*���Sd��l<?ڷTN�ATF�8�P~S�d��	�Q�֮���W��"�˶�`� ~���ɔl���Qz�a�T%ǕM�
���+͇�g��ʶڥ�=xyGo�l�:>ed�پ�s�����=�k�@r��)�D�7����|n���q�ӧ�a�)���۹�)(aOWi�t�Ơ��8yb�IY�ȏ���i�L����g�K\ȱ׼����NĚ�����\g�^n
|ȡi����o�Ӫ\/��X���a/���o�����Oe�W���
�f�V@xT6��.���C�� M�|���5<f@�c��t_����z��z�/K���vZ�$.�ڶ�u��3�%[Y�I
�(��Z	�ʲܦ7�6���b� \ũ�E4msk�	�ݨ�q�&��톾5R&�(=�h(V����c��%���k�F���(,�5�B#dn��TF�o�' Hk��wh�(��Ux&u�����:�҂9�(�߻�.Z5�4��m<SӀŖ�-d&k-Zt7�:o��%wH%�b���B3�H��o�:�#�s!Z� ���d)�l��*L�#�~3���.�]��	�?q�M:�H~����0j���]����*g�d�a�z���n'=3��P@�����rH��6�w�HN%XT�=w��4�O�Đ~�.�gbS1��`��83e�|{��#�3'(e[�g8�8�@�;t�8_M�����h�����Å�KSq/�B�w��ugR_V����cQ}�o�g��ܽ�mYՒ�շW���q!�e��P�k���g�w/�]!4�P�e#/I�C��=Ȕ0��=�5���2�yX�Mx��rZ5r��8O[�٤r�F�H�/��o#l�^x�_U��w�$,)�rg[��!if�d��~׸�Y�c��J���m�m�?�L�r��EC���+����\#���]%!r����gP�n����/X�ꧪ��d[�����꾻?v���B�?9B��%	���f��� �W[1��%�|>�kYq�������������l���՗�L@ `ӇL�Ȉ�K�S�L�#4��l�k�
v�G�xhzxF~LF��v/�w�R���قf�F��E�'���K�����M�����o	c���*�̶�\��-Ԩҹ�['�6�ە��@WݞX�iEb�!O��v��5�R5�A	��I�%o��sjBd�q����=S��O�D����(1�R�A]��.�1 �����]l�j�|I�0n����f c�\�A;�+�,��Ү�5[&܍��|	��fpw�v��ߝ��[�P�ר"�u���%uͽ�=[�ǷWz��5�β��i�����#��G��CU �hF4���R����;@�B��;�=�|.+l�����L�]"k�x���KF��K>�^@����Q�P�H�<���ӻ�ys9���Dhe.��/��T�l���Gb�!-S��Q0�,��ar6�#}����I��>��NҰԾ]�f��~����~���.)��~���s�I�������xk.1�u���v���x�����Q���3�Ժ��A�y>��p��1�C`F���腅��w
`g'L.�>�A5�R���	��a���op��L�o�ف���#��6�>Lf�m�H:�Y��?$}%��#ir(騦�ズ&��� �9�r�񬧀P��PeM���O�۞!��d9_��_|�aPY��#�s�䚮����l=K�����?�p ��m�����G����؈
Q�Z��2��#S��!���U�
CXOQK՛Y�u��>�I���@@ȶ���0��m��{f*Ϧ�߂ڍ \�}�S�/�mq��I�ے� #'�GK�MI��56s��Jsg�.�2��:ǭ�º�2u�,l��d�4�V(�] ���|m(ݏU���A@��R���4z\��GW��ƒ��#��;�*(?bY{���Y�a~�?5�.G�=�K�bXb�!U���Ǳ�O�i\Y���ğ��
�5���\p�(�@�����"V��R8����V��k��Pv&��S��D'|T��>�i�i���k'�~�}eF�;8�\�y](�Y������cO�Ei�boj1H��ț#R�o��G�@�Ʋ8��/�]�G��u�,b��^:���1�Y�̿��=�*�bl8���"1]����w1��J��)����p*�d�a�;�ч��C��5*]ĭA<g�	�&}a&LBJ�"��Vx�N�+�6�29��p���{�h�|M,�<d���޲`�]f[�I/gX�ﮧEt���"_�uX�eD��tI�h���JT���~���(�;�;6���^*��ul�Љ9.!jp%�?t�+�'���8*�&)u�?�|�@���)�$ݰ��2bOlk8�R��G� �-O�h��L:���-Ү�F��b��/Ԗ9O �q&*+5���p�8q�4������W�˼ER�^�v�%u�^��g���/TӚ"��k�PR��]�;|�<�
U��Ha�=[fT\���9s�,$lИ;$�I��P� ��F�����*g�QC'�-|����I
�E��My��V�.�2���7�h����ҸW_cwN���J�1��9�@����g��}����ЏBh�r2O�E��ˤJp#�=#O��]'�H��\�k+հ�����R��ԥ|[]^�+=�Gf:L1��d�c�9���%	d �j��C@OG�:�D��JX�*�S��=Yx���zO�Rp0��Z�3�G0+D<3�-���0��;�W��0J�f��*`���)��(��_��YoM/,��b�` �F��y2��^����-`��K���s�JI��>�8v��F���=9�_ِ��Tt�n��l�������٭���Óӽݸ����ީH���KhK��s�IN�P���I����e1v��ǽP���>+��@i��؆ !ke �v�ﳫ�+M�V�<���\���y�g��h��&9#�y5� �1������!���m�퀖�MK;�Uߤ�����bgS)�À�(p|������/+e���:_��E�T�6 �#��k<0��%�|���%[(���g\���-�FӔ301�:˪� -���(�a�Ie��Y��6=������Qn�0�a��0>�S��؊��=(+�"�'�(����h�+
���H6�T�ߠ,n�Yn�"h'thB��=H�Hc�Ɣ)��5	oX�rr�����k�[��|GC�;�q^�V�bSϻ�����;�R\0�eg��T�٨Ϸ��Y�h���.��=��N#hNT���>prL��j�$�<�����9�b��	�Nx�|9��rt�2r�%���4+r���kw��N�n�,£5�ہm/]���F-!��$
����kBT#����ŏR��o����X�2J�G<��	TY�k	��b����'rb!#��f�8��9
�9[�����'.�\�m�˴�U��~=��R�5ѡ���<�5/<W��ׯm����f&�1��;�/�Ku�?ՐR>~���=��K�߶#�Q]�Q�}>M�����KXҡE��G��/b��x��Y�q��`�_�mx'�ta���K�*�DC�2<A8�}h��%fAz��[^�4b�(�����V���#P+���t�/�6MA9<S�����W��M���U�l��妮�079���w�o�I?�a���aATB.����-ɮ�,Q*Nw�\�C�):3����	ٰ�#.�D(�h��p/_�Ύ�3�[��X���{s{$X��Y�%J[���/�eԒ�u�f���ӻP�K���CE���[�yFb.�9r�S4��{�=����$kk��WaX����3&'��)�V�D���n+c)Z��4S�����mv�{39^��C\�Q�l���#���2Z��(�`��tڄ��|�c]�M�+��b-HT�	�\V3��d�5�I�j Fs�4��IsP����R�����u�J�Dc��֗^Ʈ�1���V���H"F���pU%,�"o�������+9Y���h�Yʺ�,��L��m���]��x���a>��w ��� fe������~ �3�_]Z�#�V�C��'��w�`���hu$�6,�>�M9�;=��M�F.��͡�:/buh�|�e��Z�>Q7��J*Z�ں?��H%E�1�4�m�r`8�n;���t	,��TF�uTOE�Etھ�*��nh VaI�`�~o�����l�e6�7v\�n0�@x/�|�B�Ό	ʕ���'�jw�����橭k���?�mJ��-�]LS򓼖���R*~�Q����86Kjx5.�s
�ZT��B!t���}��Z�Agi���}E��#����b����o/`��7���R+/��+{�$��F%T%vр�*��Ͽ�=>�X�Ӥv����?��ND"��9�Pg��F�iR��JVE�=�`ʽC:]��[3M>|�I'4(9N��NIE9�|�Y�4+��1�m�"u�~@:4J,�PNu��Y�z��;@�l)����{�]ފ+2=c𑆦f?n]6v+���u;JBy��Cy�k����6�^�YD1\E���D��X������s�'�Qa~pE3��eY��]hV��UX��A��s5�
���x?n.��N�)���o�J�R�LX!� F�Z4Ɣ��K�(iWs�%y�P9��m���� ?Gfn�"�~zG\��+��Fy����|P4\Y&4��v���$mtOr]��e�guĿ,�&&�-�GYT�4˧�ڒ�BD�坘���¨,��h�u��� /���tԈc�x�@� l.��P�QK]�h6��UH:���M��'��TA#� �Ao	�6U(q�G�!�<*([ًZu_>������xo ����!X�U�m�g���By݌���G�;(;���h��1h�c�A7��3�H�Vj^^�7��&�u&���%�O[��	:�D��XJ?W��6�C_�q��0K�N��#�C��Pݧ��d�j4R)]?fc�>pR�f����w:�$���{�Sxq-t�@¬o��<�~�ol���Mp�f���i�.��<6,�*t`�l�ua(6��ԦJ�պ�E�>2�n!6��Ff��7Nl�[����}�f���o?ȃ���t� �����2��IC����/`a,oޤ��Q�Q�+D.p�ٽēm��ph�,rb��M��|.rO��E���D.,L@�|q&į�q��W7���yI�^����;N��I�&	���A��@t�L���/��a}�b�tE�]��~{8��P#�"��=�ᳵ863ژPH4Kp���s�a|m�vf�l�R��5� =�<��-��	:7d=���j�r��Q;��䮢Z8��u����@��z�b��|0Y�_��ĺ�����(Z8�4�����A��?��I&'Ȧ�X����\yP���2��=�MhC*:��+��2�7;�q���%��W���K��~
�!.��M޺ѵ �������S���v߫" Ȅ�6p�ɛ�G�(��D�V��3��:�_#��,3h�J9���[B?$|��&O>���d�U<�a���G�
��4E�w�Y��?�7�c�3����v:��:���޸;��S��l�d5�H\���ec�4c�� ��g����"_���������K@�5�;8J�1�ȗ�z�FI�PanF��E�"7}�V����I۠��JE��ƥv�"8��4��p����ǋն�������� ��v�e�*a�㙉���e�D�ά�'�DK�"�7s}d+dK���Y�C:�w�we�X/�+��P�|M���Rur��F���A4��_��\ƃ)���ed2?�1|\�3_��w�� �R��t�}t��ORQ��s3Hg���DdH���� Xڢ)���0^+�O���&�uZ$Gտ��GrSZ�U��_����2��d�8+!5��eG�/§��~R3\�B�J�r �;��@]��P i�.�A=���M�XBbTOvX_z�|5��0r rv��j.ɾ�M�Eؑ�	ʟ����3�i����s�/?ˇ���:�l��Ry�2ѐ"�tܲ;2^���'��S��A-w�y�Q,�6��(|
D!	�E<�e���1��^^� n���r�gh:�ޗzpw��ɼ���B��4 N�����.@F+k������am�y$�Kp�)6�r�q�x��W�L՛4�GO�>�3	3S��9��X)7�[}ѷ��r4�]�D+C�7��th{��7{}��#�8?Y��X��jb�2���4�i�C�9e�fO�-��ch�ZU=w�/�8K^��ŀ�h1�Ly�>{ф��h,���o*�FQa�D~�߅�,N��!%#��`���������+u�C����k�d}���gNI)+�	��	~����\2�� �T�=�ƅ���6uUI`��۪b��>[\A��g[}SB&�15�p(�c:��:8`C?6�sUl�$O;Q�ne��#*� ul>��Qpa�h&e����W3v��
����co�Ѣ��6�}�]���� fx	�,�S�r\S�f�Z��1��7��C�/�� @���O�n*?yB\U����Z�	Oӌv�ƌy���ÚЊ��9��t��t���MD'�����NW���n��)$�̲i��/I���T�=��tr����d%z�?�!���;ˍ$-��^�D����.ϕNp��У��l��hֹ�ǁ��<*
�i[��i�q03&�lI��LX�h����4�J�P�6��N� B�"���{��Ц�\9}�׵Y��fm�5tA���hU�()� �z��/��*]��S�r�{j0v,��.�h(�i3P���vͯ�8�ٹ� dc��?逨�@
pD)��� �)�������S�ϳc�����1T�v'
z8���8 �F�<���ț��ӯ��9Fn��7�=*e����m[�]K�9�A>u�~������'�H�ۇQ��E ⽩7�.������:F�i�S��[lF�u 7m50�O����X$~B�s+��O�_v�
|��WM�#x�~�;	�`�#���_�/�f-�Ɛ�*LZ��f����t�i�Y��6���)��a��{@�gֈ�zvO��[#p�s��B�{�T�g~��J�.��>������ӗ1���섏��@ko��~�@���B���d��_*>vN�2��m���"z��<���J�x,<h�h���}�XD���B�������re\|���;Wi�=�N���D�d��#.TQQ巚j���MS�ht)�Ig��	M�u%���I$���K��l�H~G�]�WbIu���H}�P(�b��
�O�+ރͶr������������`�n��*� �=`�5�$�C!�)��f��I�/,�L�@ 7>����=��{�HIS��)��DL�7���2V0����:w	Q�?t��M􉏮�^7ꚓ����\q(8G��+b�� �b���"�a`E���q�n7Ϟ��ba#p��h
9�W�m�
�i^ǒj���YT��%R�^���2�O&���N�bF�`un{�4��f*%��Z��g�'�$y������@���-_B��=㰺�ۃg���Vy��h(5滛�3>0���;;i&���(D�����?O
G�H�2�s����h��Ѽ��UV獖��1��ǟ��H��@����pT.�	M߻ݥ4`I�<��6t��#R�٪�ܴҤ@M�+Ef��u��Xz�\�|� Q�[�\]��,+���n(0zr�Zق)��Ba(Ɉhr�1MiǤšܨ�ki�P�dr��lW��R����_����=�ڎI��:[�K�X����ft���A�Z�ּ	�݊"���P

��j�&Wj����0�-�j���FK����&�s��QZ���3�5�%B��Cv]W-�=9e�ڢ_���4!R�W���mI#�/ɺ�[�n���>k7�G������A_u!ş�.���i �-�[9���nr���I�a���F�kv���Ė�E�zJ�߼��NX�C�_yڈ�������J�99�]
#�$�^]w�.��r�^��N_�h�p�f A�hw�&�}�ɎIk�M�GgP�	�zhξ��"7��	�EI���v��nl�}���V�'RL��v1�+������~�������Y�Nf۾�w��)�(֋�` ��T���
���@b-K�d�g6(_���J��WH��������J.'Ce!�?
�3�p��Ɋ8��\Ӧ��1���_Q��#ڷ}�~�[��3�.�u��n�wLA�-�)�,z3ä���_�� D�=�fd������aCi�1���9:�K�ך���nb��!?�,���LZ�[XV�n[�Y�mD������07~�e�+S�	~9b�wNqU��#H��Qk/���򱸟�#]eյP	Iس���R�eY���j��ݕ��d��G?̶�*���4�ƫ_�|غ��0�\hi�W����r�1:~\�8�3�	�"����=�M����}���0��[��1XP_?>Q�c��]
~b�'���ǅ��{����㯫�m�1�w=z�v�|(�(,���Y0�pL�۳�9���u�%��c�"�x��z���X�8����H7G}eͬ�(D���%S}�|X�9�a��o��������zA�܆u�����;d�7��.D��� L9W�R���sP�N�%� ;�%�7zKw1*Z҂΢&X���6t��f����M�|��š��$� �V����v�����ʧڇ9m�������]*|��ڣ�-��䇊-ܾ�Og��X�c�����T	1��H���=���|��Hb�E��Y|	����0FЉF��WG��aN�I��~!2+�ׯ��Z���탹lR�n�U9Kt�L%��𺻲|/G���H _���ɨN����EB���ͳ������cy[
�q�I���=���AA7�d��>�_W�����F��i���-� ;�)'��tɪ����I�H��t�`b�t���y �X!���M�Rl��,��+R�8�i��q����`�3��%Q ���@a	/l���d��j1��n��iքEUJ��a�a&b�ԁ�$�\�"���� � 6����k�;�d쨓�����\kj��ї% L��PD��cN��*�ؑ7���+��E�wY>ˣN���%�q	���ƢL,xkh_(ͺ0�U�h:7���WlTwKL�����/�E����O�.�r��B&j��?�:=ʍs�"K':>�25/$�%�_1*VgD�I�=�3��2]�Su*����M����Ǜ����r���\-�0ڗ���G��m�_�d.�W ��t�V�Tj;M��֢Q�Bn?�'p��ԟVB8�k8x�jg��xq��n	�����A���A!-�.� �`!f!�*AV;B m���~���������A��G�z(]�hL��^��:�qf�!���x�4KE>j��-6�'�nFp>��r�'q�=�ǁR�	���J⟵�gQ a3_�%Y%:_u�Ê�i."���Ө8Xd���!�C���uI����I�Н�����Y�	�2��%kk���� 0��anC`v�<�³��?5r%,���CS���z_�QN�$B�Գ�1��-7|J��U'����i��;���&wӫ��hD���)�?����[���mVJ��Ɂ+��o�I$�(��Z�%�$,�Y���V�02Had�QD}�g	[ʨ�~p�
���72'� v9�t���h?:[�U�3�"�.�r��W��6�F^����0*�2f� ǃ�Ҷ%q�2I�������' O��z��~���Ŕ�r	��w�p�A� �.\B��;(E�8�.�JGrN�����!��	}j�a:��k�s�lqp��"�'GCؓ6.�Q��t���=A�e�>���[(��ޒ�:�:r_�\�h�j���!˭&�AGQy����j����b��?w�]���A�Z�Lt테�ui�`�j�PT%��@4ր�SEUw8e���6����V�c�^[0����( �ҫU���Z��Iwp�Ļ}���-�Ȭ�߬��C`�ľ��A}`GV'���5��:�Bp�������z��.΋��XYOj%C{(�!a�Y@�Eh��9�Ų�s�~�@��	U�Z��>���H��e���O@(�\��nfB40��Y�-�d�!���r;b��a'&<~K�L �OE^��R'��NA!EgK�/��L]�z���I�γ�ƶKP!Q���Iv���:�e�����F���-����n3�j���?���[�q�N=r�m8��|:�0 ]�A��O?ca�P�"U.07Z�e����=m��*�����T�����E�)�A�C�/�n�m�[���&5�dU���g����h<�2��%o�_����r�2�}_�g��]�n<�`��:�TûQ �s"���_��q��q�·�q"Bt�l��s��i��U���Z�����(3р�Cb}͔Om�'��5�UT׹Í5�"9-��PEh<��}N���pVc-��J�Z���0�o��n�zܰG)̦���"��i2��1���t{y�f�ka4��C�|�h�I"\�:F3��^ҧ^g.�qڦ~���]䔥�#"s�bw��dM
�ؕ� ����a�4�����6G>��3j������m�����n5F{Թ
ĆFQ�#�lj,�Z��G;�j�$�q�?5J��qѣ[{���h�m�
���F_y6�F_��� _�z͸��Al2���	Y [L��CB;R<���5���c9���Y,c��u���S���|p��K��[o��#� i[�bQ{@�O�>��
�?�Z�L[ڠ,:U`t����!nmH7�O���:Ϯ��D�ƈWi�|�Y8��*k}�	i8�G�L��&�|0��K�.'+a1i)��P��AB�33�ɪPs �ʨ���
|�{��X� ���V@�4x8�b���u��Z��!}��F�`�{*���SS�GJ������Z�V�e���(4�$�(/�fWu����3�za��h�� \��)�nk������	-�G	ī(a1,2�G�>�?8�aQ+~�� ��	�.G��������P.C��%��C  ��lb���J�6�g�,ٳZ���1���r����I�ؙ.ak��3{���\G�!�ǝ�'��h��v��/P�4�ߜ��h���,���%�����K�"YQ�������T�R��X��F����wy-(C���-[��U'�t(�h|��>�w�}t#P��}����(-�R73�T%��_�pv���j�D�Y��l�S�R��=����U~���B�ꥁG�������
&[� ����=M�7���%�T��PXsT�pEȐ���N-N"h�t�n����1�p�9N�m_��W/Vo	�!�Pf�b�uzc�8����0u��gh�# Uҙ���KŹ6���1PA��K��=\n�ڇW�a�ypk\
�	�J�:I-E�m
 �8�:�W�K�"��f?����Zf�+ek���ƅ�[�Y xJ��������Cx�	i��%��;���ĨP�f�
�u�i[H,�� !%M�Kf7h���T��k DM>56lb'�ɠ� 5jG����6�T�ݖ�&UM�)��W��[[�v��J^��sL��"�������eD#J� y�3>-ߝcD	�A�/
/?��ixV�mb�s<Uݏ�xP�7$5̯�:E���-kARz7}?Zxzq����wg:ӱԋ<~�6�m
�����P�����]�iU�ST {�Ǎ�S�)#���Nm�O�E.z��7�x�/o[!>�Oy�g}� 1&�)��͊t�9r�%{İ�Z]|��~�]a-"�{n�**RVS=[���=�u� ��=��D�N��#8b��on ���m��ҒW'�v�į֖�'���2!J��Y{'<EvL��*���-DvP#~c�E�.�k���JC�gZ@h;g(g�`�BJ<.��Rd�z:M��}���P'���#,�HB唶�ٷ�5V��u�N�vH���	|���Ӈ /~b%�
9u�+T���+��(�Ҡe��7�*P��U4M��Q>��U\U���B�롐đ�*h!��U���R=l4���=��'� 9@<N���V��r̭3���-GJnл�u(�Me�5�r��������W���o��X'SNy�i�\Un;���ox`䠡��q{����RyM�����xc"S΃r�w�E���[e���Հ�௅z�ps�k̾WT�v��?.�p�x�Z�TġA]Q�Ɏ⍏U�uU(��%f<V�3��s��@I~[��kӵP�^���~��X��;o���XA=q9��W��	3(��O�0F�Iwӊ�7����pה�3��A��_�#o0�I�El�?���^EH"��$W�^W5BI��.��׌�!xX']�O@<rK��=ѥI�O�ң������@l�1��*4�B��F�h�~�m�w���j*x�#u1���,)t���hF��7q�m	Y�1ɝ�oE�Dc8eA��)\B~̹%2:�ೂ+�S)A�/��������,�bN�≇3^�k�:ɖ����u�HhB��$Q"��>��d�Đ���B�S*�����s�qP �N��
@Q�N��ELry[��
�#�zb^`�T�����ɻۻ&�A�mQXg0�EBfo�f}`��
ɯw�^Y�������.�K���w�׏���I0�(<�5��̭�����¬���D`5d�o��`�l�p}�j)����y/�q�F�Ԋ�Z��K�g�]Db�qڤ���� �J�-t,�)Gıɐ���mƝ���tq�n�f���+�?(i�U<%�mhM�Z��?#���d��������H]J}$�o5�/@kt-% ϑ���h��Ql��
;-�h�v�!���bǦ@��5;t�cT=�Kp���H�$奭�ťǄ��M͓Dt59�h%�ٿ��Ao Y�RCo)J�R`ם�(��=���������Ny8��9��rI��i~�M�,�p����m�hr�x)�w�ikG��G#�l�Y�v;��;>���vq�
[~�m�Hv�_7K�X�ُKOB~�l���i���w5߱w`甭j�t쯺xB� z�6hJ�R��ײ�,�E�%��񟍝�	�$�'%~6k�pRo�&/
��Ymk�3[�!n�q߂��[� *�"��3s���sn`�{=�Nh�G��A�����4��&����O��"q!�؄C�����Y��^_�>�����5O��Pr'n�@E�⍞ۦ�jEJ�4,��L��I]l�a��@m������.݄��'��i7j�"�h�5H�)r(t���z�8$]����xq���D�0�8�QV��T�pXۣ�Yɗ�W�wH9`�@k5��аD��)��x;�	��T��0{a���oG~Z���d����r���p��Ί�����Ȁ��&m�Ph���84i �M�a��l�צG���7Ć��0�nڅ	��U�� 0R�m9��(�0��奇��L֛�z EJ�I�y�g��%RC��$
�xj�__7���=#�n�@��\8/� ^�hTة4|4l2$�*�PTd��{ܓ���<U�o���r:���.Ȕ+8��ߦ��a+-ލ��4-�[7����@k
;>K��|���L72M�Fv���~���2aD����%9�t�g��͔�IHK�PiC�"��G�OV �Ұ������Z�|X��VG��JNK`�{����0Ŀ�XV�밬�j��C]fcM�B�a��JA�ŋ����ʻRNR���BBT�� �9;��G �]k�PT9q��������k��f�iH��EgL�z[�����o)}�1�1!��)��B��n��e��H��Dh(b�~��v-�ͦ�ٲ
�"(,S{ك��7^מE��s���օVJƼ��"�F�Ӥ5_~ ��֫7��ǕL.����T�ha��#p�����8�0J!�F*1��ظ��5�Z��g���G��l=�U���voH��>{��:0��9ۤc��A ��0BZUuAl*��򚯗xg9.Fb��� xq�TI�J��T�XM���4�ޠ��N�V�,p�6���hќ=�)��j��l�fy���Ǫ�����!l9�o�O�|C��l��e�@�9E�=��΢X$$$�T�z���U$|v�#ׇ7�W�j��v_�Z`<#�́�NG%g������
e�@�������c�"Y=��-ު��c��¢Rc��%W�9�;�o}��Z���|t=���\4���9��:V��$���F�����(2�ήhO�:$�9��g�����:gQ������P�2�$�t_MKY��6�'3h/D��q4�B�t�Bb*f',����\tl�V����6�ݡ��:�jϊm��s?v�x�� Gs���_��S[��1Bd�
��bP�t9 �%� �HVu����+_ϳ��t�H�ә�Z(5�Yr$���C�<Gf��su�P!������Lߝ�*L=Ɯ*�]7j�e�I1��u������5t�Z'F!Dr���[����'��˫�pL	�V���[N��B��̨�=Q��N���Z�-bTW{O���#0��M�OO=���#�i'���v?���<T\�Z�
�w�1�w��&���/���������O��|�˿����sO����#�]�2h�?%-ܒ���`���K u�\t
Z=������w���4��Y%�E
׏�%�?s��J���oe���ƣ/i�)�|g�0��JK3����`��o���c���fl'7ɮ�B�
'a���x7�k���]O?�GZ�_4E����I���3�#����XX!��Mޣ8�p��F2(5'�"8	��_܊?�G���7��_�6H}]���=;Oi�Xn�kA�ڿ�IK�w��4�6�	 �����{���.�+���-NNK{���u�^J��N���ͬP���4�������i6�3U.���H�ޟ�\L�Iq��'_/����.���/̉�:�����v�c��w{���iZ�:;kbs�L�'C�C<�%i
b8�y����J~ju�U ��gwL�4)u��oN�
q��I䲤�!���`z4	�C�	����Z�!� (�ï�S6F��ɘ*9��J\��폓CˣcDc_{yJR�&T"�~:�����*=���Q.�y7�c{�։�gy�X9��� 4�}�]7i�Kቤ�؟ e�l~�)sPb��&%x�\䬱b�~��a��)�0|̈́�'C�7�y�·�]�q�D���:��J����?4�|��^��u��׿�����[�E[�j��j�j(�و�2$�j�H�ǔ���BO�N�ei��j	A��q �0���^M����t��J�.P���y�G�6pe]��u pw{܁�g�qU=�g���s7�P�
��|ɭ��/U�Y亝�$����L�۳������W[������Bi&��A,�0Y�%�;rzR��������?d��� �	ڿ��60I�},�]�]Y��&��2Q����vB��f�����4��:�_8X���'l��v
O�Uc��֗���p�g��
~���~����Y#|<"���6@.5��q|3�'Y�f�R�{A��u	��=�6	���T�����1��z���D��K��ysQ9{�dw�<[���&7�d7�����&Tu� �g��Vړp�e��h�{L��ʘhNt�z:��<�%o���'�_���PQ��D����,!j���I��iZɑ>�̕�M�O��@?���q�G���c��S<6瞒�0���DR��/~�'NK��g��f-��
����w�8���>6����Ԝ����[�Q��J����S�A2Po�L��T*1>wj�>���.�Z^�vb�P�UmK�&pxH�t$E08�©���?�� ��"��4������G��W_�� ���!�*x/Q*���ت�^�N6h�a�TH|
Qq�W�5���y�����s��� �"�#��ЇS[��ʩ+XpOM�R����e���dzD{&w �m�T�y��"4t?��E�0<9���{*Q[��S�����Z��;������0���zP���^��?&�N�v~K��@`�3����@ۋ����u
�ꏌh\�%a�X���Ocz�I�D=�.��4�8�L�+.[-�r�ú�i�tZ�N�B�3E�2����Tu��}Yۆ���1�w�y�����m�<�&��i7p��S�1�e���~\#\i�&�Z90-��jD Lw�C��Zw�4��Ϯr��N�e��y?uJ,r]�_ܟ��(���W�x׾@n\�.{�I�i�U���A��BP����R��e�1�,=�k����~��Dp��_�uԜ}QT���c��M�f�,KW���(��/����>��I;�}�Gd��P=�t�ʀ�r�j������ز��1��A��7p�p�*�f��� 1?d����W�d��AÓ�:&�X�hp��5)?�'�aXeM��\�j��|�l.�(��2���k�aO�� ��E)|�Aȧ&6C�tU�Ɗ�z�z����8�nݫN�j�!%x1m\�a����y�:(��L������;�yrdɺu�MŦ034��u�RZ1�9���L�A�GO�z,Cr�L�҅���B˺�J���E�&�0JMZ�iJ���~��	fȗh�F<�S��B%��4EL�:8wagaɍ>}�J�NMF��OtP�.��pvΝ$go���8��T�K�2J���:�Y4^�28Lk�[K�fD` ��3/��ۺ� �B��ce�nt�JQ]H׏^\�e%��������_`�y��{��mcoaDwE����i�\3�i\E�ۈ�#�����f�yaY4�x���٩M�-w�L뗰�T3S~l|O��=sL�%3G RPa��5]p^�\ :���?3st,)��!aH.���8(3z���N^���q�5�O<W�k�GU{�4?]}-��[����¸���=+~yk&q�"�o��s�l�6b`��K�����bMX��p&˭�����c1� #�����q�5g�u3DF�o�қ�k(�yt({&�n0�|U�92-��׭W�:=Ӣa���>-��W����S��Y2X	|	Ό�ĳ��+�8�N�ߝ���p����j��
m�Tڄ5��W_��@J\�rg"Hv��EJ�!�q���9���?A�`RT�f	�?�p|��n�kb =��ߋ�N����P�L;�*7Fo��b�Z֭Z�gl���ԯa��)Yn�+�������KC]�9/�v>>|݈��[[p�K36@�2�-a��	�#(K�eKŋZ���[/�z�ޘB��A[O*'|@��į��cѕ�$��ޅ�k�2,�,m�|��m�/��=��ۤ�(5,�"!p��\Z��#�#�^_���k�4��d��}n%��7c���ƞ��W����lU��N�X���T֔:~w���\���`�4:��9A��9��ö��<�9l��m�4-�7z]����;ˣz��4�ʺ�j�d7 j���k�Ti�fD𳳸WPx~?R��&pt�����r������瑶���)�N���L�#�a�4�p��tP��o%�N*a�0 Nm�L��	4iF���O��2��Ó�X��d�n��T�r�c�I�9b�r�'�@,�R�8՗��?��Y�j���h�<6�Q�Gn��Xv�e�
8?�ի��T��|�x =�����K Q��X�a�v�J�b6o�e%P�+��M��D����W(L��P��
�vRl�l���˹,�N�6���}�7X���k�Ζ?n.B�0�ބ1�o@�U���ߨ�Z�P��}�ރ���cta����\�M.X�P�^;;{NQ�h)�����9�ʧ�J��O0.{�����Wu�z]l���|Ӌ�Z�d���J�4�K>�jKDؾ`}�����a�}�@��H��$��޶&�d�NH��I�����O��\�8�0��� ��)���Ю�~Ϻ$}F�e��`쯗n��%�G7.$�8����0#xɎH����YJu���k�����,�+nEO90�+h�z���O�Qh�ܯ�ЫAc(��:g��>h�%l;�.�yB�M�>�#�hO�����K�_Gf�]������d+�Ԧ�j���bz��.bn4�<�� ��A+̘;��̢V��4���IuA[�sik�B��^�c���Ԙ���K�f�-5�z���3���t��Ue�)L���dۣ�o�آ< }��?�ɦL��⩸b�����z�$�l�.>�ֶ�]��H!�U'14��j����O�`(y�&��p�R�z�ܛn�#k�a��t~�o;��|$ցzΜ��#dg��9s�h�Ф�]�<U}�S�~nD�c0����f�JN�~�e����Ցb�c3���������D���9P!��r��}���h�x�*pv�7�l�?]���[1D	�v���3��%ԁ x>a�j�'6�����a�����,0k�����2��c�s�}[��΍���͵���)S�v��y��c�DŃ����H�!%:y�P@�o��?�eՅ����&$`:r}�m��ɏ�����h&+1�~��i�l�q|�F+�/sM�|�	�Ҭ�K�!/}��?��Hop�*L��8G%9ov�2� ��e�����	By�^-�i�},o�O��h:�Vf;<�(g N��!���-�P"�<h�5}�ܚ崑<SP:c�&�"|��e��'W ����P�������HjԉV~���mi��cџI���pi#U�7�$!0	�����(X���p��"Z�r���B�o8Y13�$z�A���J4Q�HURD!�Y�:j�;�*C��{ Ei�ʸ8 ��c�J[s#���z d2,�i�l"�|�%�a��x�Ϗ�-i�Gr"2����vM���ӭf�\�>N����," |[�YZ�7K��%6~m۟S��`�"�u���^0Q�	��2I.�L�"F�<18~&>y"��t�>���|�����{��4S��$��9SWL�7�k}���Gb 0�v�%H.Lk��j2� ���D�K�WO�Wɷ�o|,�ߠΕ��${|�Ԕu�<���Ƈܻ�C��J�̟-u�2L���]�akYϚ�s($�8hn���/�t�r��0Z�eӫ���� ��+q������y֫4*Z��(�Nh��]i�6Iy�ȭ�[D���������S��csx��ع���G�Ų=o�@r⦊ ?�`$����a�<$���6^�-��(�ZJ���"�N���7�ˤMʯ�4����Lh���w
��=����kTdW_����}�����U�,V3D�N8Fv�㑩�:��+d����aG��M�����rK���t����ʃ
4���qH�g�㝳��t���6�B��"t�n�庖:�bf�))~���p�4�u��e@�N�,JG������?5J�"f�7�Ls����fmz�X�����v 9��7��N8�\T!�g�Qʪ�-���������w�6��]�d�A��������:ë��8CJ�sn�=��Iz�ɕD�U�!��Zy��X�ɶk!�j�A�A�����AD�w�0�2�>�y�΋��nz�>�6	v�=���;���i��R�J�G*.:�v�L|�_k�qA��Ny���=�Y�>����$�#�DYU�����j/����G:�zX3��'��\ka���?!y�?��CX���#��[MA��g^{p��ӎT?=!�Ju*���\���ݺ\z9�hX� ��s��d ?��\�ǜ��.�[�I:�v�h!%JrO%���9D�M�C��-�İ��)��Ǘf�8�`$y��D��3��>H���\њ�!���e]������}qm'wO�����=�j:-�@%{e���� �/w�Q���H;����:m���)��7�%�\�����9@�w�;6L��)$5������6�����8������J���	Ӷ���X�.��[����.?��ؒV��;�L����NO���Y�![B�I6���6�����p��ɖ�Z�Kc��������tӊ8?�����F�F6Դ�0��B>��ˠbA'(��H��M\������;�	4&���h=�_b���"�r��q�Y��䑬���qq��>�._7�~�Z|l(l�L�q){��)p�Ee�d��+�뽚s�6� 9Q�d��e����{����8|��A�Z_����F
�Dm2���cy?�2|;_=�	�-[�^0v7~�Y`m�F��.�	��`���p�!nފ�<\g��1^���c$��`ތ���a8�
�O�9��(����;pЍg���Z�.�X�JW�d����e�{D�G#��e�.~265a�d�j$��X濽��x�z'(0���5qLģ�7��7F�c�����<u�c׍�j;�	��ռ���7��W\�5��d���Ҧe�O�U,�Nx��<�X��x�o����_ +��ә8�jL�p� Y�H�ڄ6WZO��y�n�(��{�TY�yp>/�t��U����x�:��?�95��u�x������{�V)�}B�ͽU+�7*3���w�9��;,K'��J5܆��ۤc���p�N�n=������BxwP�h���a�5i5T��[I��t���}��5S؂�z��C�i{�	�N��~�k�'��UC�O�K�������)�:I��oD�:���em��/���	?Ob�Jx;P��"¶ n����r~����
�M�Hy��1���C!��@�rr	p�ģ��.�QǎQ�נ������-I,u[��˄��I��B��O������6���@F�G����N�.쪕�4�w�1�_���s� ��Mù$l���q�[+�I�;������MLؔȚۼ*�9<B�o�i�z����P%m���&	�<%���w�x�;���=;O)-X��G=m��P�1V��?�[����|sK}�������΢�|��m̛��H�`ȫ�
���_�����5@�TX�����H�Kx��%4nُɓ�ڴ'�3z2	�:�\��o`n��(T ���ف1A740�� L@ ����=�/�9^ ��ז.�a�I[�&K5V���ZV�������,�fj����A�B���ǐ�-vn@��ZYZ�>�c?�J�?A����%�4�;����_�sPg�l!�i����ʹ��Fq� /�����@*���N��D �X�F��kR/�wR\5�o�@����Qꕐ�'�}b��yH�l"z��ɞ��4��3��Ga%��Z#���G�ۻJ���(�7�I��)9����dɻ�^����5� K�!⓸RR�ax��ؿ_�4ķ~PN�6�n�(�W�o�	}nJO$������z�E�����X�e�x��-�mr6}�J��m,��y�F�b`.��;��Tc�9�|נ�4 �˩!���&���HdU���l����S:_*$g�I*�����y�y���=A��� 襣5�uQ ���#���)th��Hz�QcKw\�"���*W��,h#���H��Dސr��x�ۂ
��L���y�n<�gDa��#'d|4�W��y�YU`I���	�?9�Nz���U�%��`eF��U(���z�Ue1��"dqZ	�P�(�Ԥ(f��"�[�>� ��k�}v������c"�{�W��m0�5oΝs�e����Dx~zU]L�����BӬ�֖ň��Ǻay�ጱ�[��ώNX���<0�$;]�� a3ib�+�{�uB?h4������̐�zOШt�H�i9<f�XI��,$M@�̘c��U���+eŴs�,Ya��Ŗ29:�ҿ�wK�T���L�8$N|[��"��2p@A�jR��àzo��5�M���hn�.�-C7�z��q�&&�R��T ����\����_���$��  ��h6�5
*]g"橂he}Rv,rh�d�K%(޴�3�9���8��]d������k� V�bH��X��;]�C�$�9^.�Ŭhv�i�#���e�t8�h2�.�-z~�t�k��y"xc���w��s�}ވ�%Wt��� R"��/�7��� ��dܦI�`��������"�c����MZ�^e�qo�6�G$9��O�]�La۾K��
,���\�x~��H�@/3w30|#Q��^h
�����]�℣�ʼ�9�o�Q����]`���i�����X	f0g`�:�k&A;܉��ul۶c��8@�w�g��x�j��}~�V�6丑�����z�E-�/�4o�ڪ���O�����fD>jC�>����n}yKU}��#x���Cې���K��.�%�{9��ߵ�d'��Ӽ�A�Sktz��ӵ�1�������Zg3v��$�Ǜ�� [��n���Z*���zR�������u�P���V�a��j�e�m��ϕ�s��X��K`��|b��Qf2C�Z%�!I	�͕-�u>)�p�6i9���2���#���2zZBn�g��u�ou#2��^�+#'���BD Ӛp
{*��WGa�i���u8�\��h`u���JXE#
h��"~I
�H��ռ�u3��}k4V���ǐ�N�e��^K��4�<>�F��p#��z��/UNұeEt��:���^��QH�$�F{�#��G��:��r��fT�x����P�scC�s;t C8ǎn!o��3J�B;��";��߅�� ��\�N��?�c跰�
���z���O&�d,_0�18�6
���=T��P�o��3�ӫ��Q����n���FM�K���@�+r���S���1a��c�f=��ٌ��(���B�G���|'mҷ.-��k��<I���\��v0��y����W�P�nN�b�<��_{Ea~�\�3�6k�6�G�
m�m��=�fR}N��b�A@���k��'�}xz�������o�RF��hD�����b�a���͹�I]��"$����Rlǣ/��c�]v�5%��t�	��팽p�~�F�{҈<�jQ�s�������h;�N�y��sT~&��< �*Q��0��`j4�
�f���T�����w�!�2Ǥ7����7�>�Inu��Y�#9 �/��`u���>(p��c0��C&J��P�w�r%�˗V�Ü|hu?�z4	��d{��L�0���	\D� �ݨ]Y�m(�
4aL{��~ce7��a�M���ϝ�ī�s���L���<x�kN���sơ!�"��7�x�M�m+��E,D��O��>��J���0��dy��t�����Sx'����P�p(F�!�Yla,R��'.�����)�G�������H���c'����'�"q��i#k�ngT�|Y6XaL|���k(�ƌ����R��]��.��!���ƭy��(�(��x���ڷ�6O�g����ä���b��1�D)�܆�e�� ��JƑ���ўk���KЃ��Bc�)�dg�������H������g)��K�g�6)�eD��[�-�;l��s�a���3�k��׹�.І��h�2NR'My���k��6s\r��ְ:��m:�W2а�a��I^=�Yi�N�1�4۾#�Q?���@
BHy��MF��=/! ���;و�?P(g�mpH  �I�v�l�?���e��Ɏ�.id,�_�|;}�?�U������#n�(1) n|��H��,ƈdFp��O&0N������D+v �F�l?W�7Y��f6���zQ��:���J�!�B/x`�g
�ps�7L�El���s�y��~�z7� h�w��F�m�	a)b�xSY�)E?߰O&ey`}a��E[D�TN?�A)*���M�����B�����j�@T�{��~����E��lc5������Uf���I�g����4	��Tyʸ�&�SФ���ކ�X�֤h� 9r��إU�"��;����no��c>�(y�F�������(��t� �)2�DYӳ1���a���@��_�W�E�j���_�0IK�.t�X�x�[����|��=���ū]��� ���0H{�.�}�M�i{Y��≄SY�V�� MmY�W.+��0g�7	ng�p�?>-�0�HJ�7<��ە�d��J�<�4�(���Q�]�O�$��Mi�/p��#&�C1���;R\yU��W�@��
Bm�La���0p5;��g�=�TXā,�%qF�� =�����w��Z�Wł�k����C��ׯ��}�5i���S��l!��N��saB��'Qg�/2%�C�z�m��Q��}�SM�p��|���y�7�,B�*u��K�7���A� %�����c$}qq*b��$)*f��.��5"��a������kns�Ln�5����As�M�x��7&v���	�0<T��dg|�oP�;hP�a��=PD�]Š�_WTP��l�.!�3�
��ׄN�>b�=I�M-�����5�~G7�Y���\�a_�>�нلZ���Ն��N`��4� ����l��7���CU.����]GC~ ���e��\w�JD���w	��	f��쪖�sv�E��(�H��N���a��o�i.���ͧ�����J|����|S���PNG� ��MC��Jt�ȇ`e1$U�hhz4E�* `�\(�M�9s�u�����kZ�P���@�8��� ��Ș\(�i�2�1��e�od�Or�s�L�t�o���݌m-�uVX�>;#J�}�g�3>���7���T�X�|�E*�ɪ���U\����#Y��8K��Vrݍ����C͑Ȕ���@ĺ����bu�x���ă��1O������/*�+;�@ɒ�TClA���Zy�B�39D�l�F����4ta�=��n�
ZyS�w!E��J�>$ȃ�`�o 07I߬w}B��K�@E-�hR�[��XS�6�dqěM��|��3�'<�,'2+�rL^��3��<����hm=�	2���z�i���s������ر��h^#r� ��ݘO�Ȭ����wXȮ��N< [}i�����]��+��+��i��3ed�wI����S��ěц��!��D��C8�qa��)�6.��������<�ǣ��qSs�F$r�x�{�h��ɍ�z����:X���&�˙���.�����ێ��'��;tN�0n^Q���CPGZ�S��ݼ��%�^�I)bd�Z�p� ��wC .�'i.i�3It�e�nuZ �8���l
��g{��g$�9ɕڊ!�L!Q	1>��g�n�(���N<��4�]
g��ߕ����_�7E6D�/��?�0��FY�����cO贻i���,���CF4;罝1���h)/ �N~���Xz̠qG$A�@K8\#��g��{Ni�	�r�k�l�P|ߖ����D+�>L��c6�ewfFGX�g���QB5&�MѦ����@O��U�h~K_IyF�Ћ���{�[GjL`.5��d�p��৽9|̠�7�{�?�)�ӂ �EK@���}B���U�yy�5��j� O!Յ���2�P��cfr�4�4k����9��C�㖯�;��E�ی=�:� ����`��z�N�E}�k��i2s����2z�Ul���U���
�Ȯ�T���	����瘰��?����U��"8�L��	A�%���	G�2��J�&)}�'����F�.f�實?v�8d�^|�Q��&o�"�����0齁���8�'4eϾg�ߔW�&�X��y��þ����j�=kң����-0�i���)l�Ãs:�W��ď��V9DdeH�k<ut��
ÇC��n	��,�Ц�H���^0��mL�$�̷j��x�2�>�\�^_>���{�UP��vF?�B.����a� 	��V� ʫ�$�w�7�E01N��wG�Kd���@@�E�$�=�1�.���-&-�)��լ�kN~h=	��!���2�Z���(X����#+N������oף�X	��7:����!�2d�R�u���ph��~ �YZ��'�/;�����1�8�zfj����K9�o��4��nd�	��o�#�&�˜Qf�q/���,�ld�;M�N�?�����M��/�y�֎��@�3���V��#�!CU`v;C�C�!$YM���S=����#װ��aj] #��ḟ�E4�x����@N@�ӕ�X�9W�F�l�+7�ͣ�`hT�ضA�� o��e��^j����y+'�!����>�z�KRr�甀�y�X?����XwBܝ��n$������P��"6���;u^χm���b����{����q�\���T>���
� R�ˢ�'�w���Pa�چZD]g�w3�rn��,��?��\٘�f�|��0HJ�V,5��	���T�dХ"�K��N��=&h�:w�H��7�mQ�l�zZ����.g�W'U�e©�CZ\���%Yi�͜+RH�n�+W�S6�{���w�4@V������iFt���2�׋Ζ�p�È�$���R) ��&pY�}]oM������XM7��%lD�V�R��7S��U�(�;��A;�"�}��XB��RM�A��?���H-<���n���΅������L����1 :�����u��z�n�/�����i�M��+��F?B\�?��E�������;���)��)���=�YϵS��gC�c�T�뎽��+J=�Y����J[�XZ�E�Hgdͥk�d ���=�x<�%<�ȁ�i׎��S�G���`�[�9	��؟_	��!��Po��4`Q�+�%��m��c�ŇW�FD��A�_V$\���_���z�Uw�4�*��-�b_əOsT��	Z�~�w�K��f�sXy��j���
L��=��������pF�b;��T��p5j�WK�ki�ǣ�o�%n&"�:���u��i����^��1�,�k{ңٟ�����<,���ϻ�v&�Z�����ː���CRH��6Cor�Mɉ�VKͭ� �_�J^��4�f�7�/������ͦ����U㷬��%�>F7�%�ZG��c�����AK��1���%�-8&w�l����V<�1�<Y_%��\����M��ِ����8�O��0̋��JB�д6�-�xP�Qk|4ˀj�����-��}&�w�,ح@�1
<JSt�R?_1"��	��V&ïQ������?���ڏ �X��&��Ok�i��K4�r�2K��J2K(�c!j���3�;S�/ú@6��;����Ɣ�X�-z}�	��j��|c��A�-�0��f$�W��� ".[����F��9I衩�r2���Z���<2;$1*P��f�5#�����o�*����{V~���b��?�QҼXeEýu�`����ݘ�����V0�Y o�ޱ|C�!b���UX��n_�����v�_H�<7Ͽ�[���E8�Ary���E4e��!�s�������S?6��؋��sw��*�(��Sa!��kci��S9!��K�Ţ���Z�����p�&�����<��&Φ,�B�YZ�&�?���j2w$X`Zީ30`י�k�K?��̐��+��knj�6���3Tʽ�C.uQ!�g3 j%+�rh�2m(�&��'D���Gu�=��Ф�1��P�ﶫ�����/�J+�0#���oi�5lS�"a�z[C8�O^N�_�O+�X�$��OW� @	�w��2d>����#����jQ��`5�T��%�}$�zc���[���;W��g5k	��,d#Ô���lV��������&ki�i��j�Z��@���APN���1)���\<�wT�y��5S<ɏZ��V}�Jz�#�� ��{��!�Cm������7O�[�
F��g����^�0G�H���oR�7u�8:��L@���z�#~�S�Ĥ���Ud���VX�,!�(t���T"P�8$��l��
U�K�����MJa�C�
���K@-)"��H��2�L�]f-ٛm=|��M�(TR��[���˕u���I��ˈ]Y$��LX*&���l�粜��X��S��o�r==�g�YI���ڊؼ%�Y0�r��J�s_�a�&�Ñi��������!����{VwI��&�Rӛ-��'�,� ��/+�n̴!rEsh`�VČQ5��>�¸���rb��EO�d��Q������FTa/򰕲i��:W��6�/��\D�RP�x)0X�*��>�	q�����Z��@'n���[M����[O*�Y4���=��FG��&����)c�9���p�l+q�BQ��dU��ԟ��G��H(8v�1�&T�A[P`J�c~��ٳ�XJ�C���W�K���pL�Ivv�F)��u��1�\�q�ى�2�k���P��������k�«.�ڋf��wy��^h�M��}� '�ȵ
��K�����H�:��K/^���;!�1�1 �R�ߟ���}/��B&��2�P���YE�:)�4.�`i]tt�N�g�cV������I@n�\ҡN�1��'��L�����F	�Ey���yY؂�T^��fNj~ ��ts؎3�(��SXn"u�/~ь���\�앾���vְ���4���ˌ�Gn�B��@��X{2�z�6�
��EI
G��a���������%~���=$����HOfɧY^!!�D�QEb毡k �"$A���_7;��r����or�"-W�п��
!�f���N"G]�(<S��GЎs���&�q܇�/~W(T���KW�$+�o�2��V�?�D�Ċcߓ�����}g|L��J�ԁ��ݶYZ���8Q�M�����mlE�����G���_��{vd��������H)ݸy�h�掑�c��
^�+���D �"���w��Q����;���v_���YN�:�13cZ�6fH��+s��2���xQ{�E"���L�*8ju�=	Ƙ��t]��{nhS�wm�����S���
����u�|�!����F��;V���`��qt�j�Ki��BB�p�4
�.C���Ex�1J�$������ �̩�k	���5{��z�8����I1�*	ʅ4���玸)�,�i=�@B�~>'�M�n['^�(럌�{��-��}h��!M��V�a�>|�Aɤ`��li�61�z�Y�ߟ1��k`"��wd<��~K����<�=������+�>���ȥ�c����	�������h+���=��ş�k�hu<�l\��%U�ƪr�B`��Q��&r�GDp#s��
!$TR�;P����ýD''�9��a�\���e�ɕ`L46��S(��1Ϟ��O�zO�ն������tq�6m1�y%�)�N,Q��g'�P^M��@��u���,+��1�,����aІ���}tc7��������q�%�c���2�ț�<'O���6�9N�L�?��e$�o1Һa��~�q|]ȅԷ��m�=p}u��Ε�fR��k*id@)+�_+����?Z�8����vfZZ$���.=&k��~<o���t! ��=l5��իlT�'�z��T�s�:ze��@�YZ�E���*"L����$����t���x+����?*��fZ��ZU���W�0+̃��B�bZ�&,�>��i'ۓ��-�aYp���#�-%����dk����O���\�l�8y/�kl��9��'!��n�+�4,�Ͼ�/n4�zBƞ��"r����6�"뜨w\Y����� /J�\|�̈����0��%�jq~�|�:>X�o��N�M���冶g�����Ѐ}�v��<�G������`HX0��v�[9�CJ��*��x��4�
ю�~�׻,+b[�?J����*��W����O�q���8� &~��nl�Ғ�Z��YɑQ09�4���=�׮��<���ya������HP(<6n��s��t��( �2N����<	�zV�w�M�ٲY���ƣt���4%�D�z	Ԏ������2E�c��	/V%�L�
��̢qw�|����? ���N���T$��ʪ���{L=s��!*[`��Ms"�-h�yNĔzEe5��N������߬ζ���[�_^p�ȕP��iO���y����B���3���X�%�ph�!��ᢘR �S�c�"���T�����ۚ
�oO!T6�&��xؑ�X��ũ�C�%?*
U,ܡa�{���װd
??���rՆ���[c[���5T�����g%�����֐���=;�ǩ�|���g���g��IS���u���[������!����v�3r��ȵ��
E5)�p�]zɑ^�jGW	�T �)��`[ M�����k>̹���Vc>�L`�x��y~h���ՙ�_ ��V��]��	&g[�?�������v_��aN����Ҭ�W���1m�p�\�zpM>H�Ɣ5-?�F���Sջ7�E��6x�N�U���-~�/���晢
d�Բx@̽�w��c�K>��[� �L�d��]�a w��>!�/LR �ݿ_���T8���������⊯���&F�
$&���Rdv�'P �}U�qʲ>���t\��B�����I�I�#�Q-��4s���Ϥ�\Spƫ��	H��i���;⃊���-��u��̆��X�>�+��q��MI�A����j���m憙�Hh���������3�N/�@O�nK'��~D� �p%�J����6iI
DpàA�����;�n�Ջ��^n4�8�
��ӽC���հ�>�Ȕcq��!&�F`��'����!�l<�����޿�t���G���vr��0q���$|�L�e��3!�X�?��6�f��I[���l\cc�p��0��	��#o&yΛAڒ8`v��h�	S�d�Ŝ��u���}��f�]��FryN@��8~J?`?E��/�Q �3�w���x�J�%.�O=��{�dҸ|��=����hW%�a��k��x�*R��_�i7ڻ�Pa�ӭ8H��ٛ���M������.�|�#��٠�j���;����V�!��Ns�j��z~�[(y֯v��v�}��a��{�8�s��S�/��v�Qe%�f������M�3H�¼�ܷ��4²���I�}lҺ����r��a:�j����53�aNY���RV��kP.�k��K�i:��{m�LR����@�Z�q˜���9k녧�ƴ�s�o�!�$��4��V���J�Ya��E�{�hx��!-��Ѵ����z�2�Dl�S�3��IXƗ��`�ȁ�z�(�,n�V��Q�Ɩ�I�Ǎ/�0��݈�x�x'�<�AAb	��O��[c�E8։\�o�^��y���d�8p�m[eã5x^G���s��ۃ0��Ll������7!�3���3��r0c=m���Q[x�̀r� ������lCa�V��O��%���� �G���o=�n�.: P�.c�
u�W�*������_�oߪ����@�5/Z��U܍�N�a2Yg���-2u$l<�b	J)�d�HQ��q�1�7��W���{��$ �ZА��e�MK��s����ٞs��݊Uqΐ�-�����9����M-�9_uP�9��Җ!\\̐�ל�(�v�n�e�[+x�nX�Z������|�a]�4�>�������
@�,�lk�1M`����r�A�	<��*�Fⰲ�L�.Wg[w��9���t�F���^�(/\ ����z=�&Oe�$\�����>�߱*�+�_a�֋[��\ӊ4mɎ�(笳[�\�A/Jn�+v����Ys�b&�e6�gB���3�ݰ�e��*;q���[�����C����p�ln� ��rQx��Ut禼	�?񽉶�O��_�|I��V���BzN�2��$C�[ɞ[��Ma���=9�C�o�a���w<�*���a�s��jJ�.��\r>��>�+p�#M�����n��U��P{�t�M%��X�lG���H�t
}�>og��C������t���+�QɞJ]�^c�?�����(m����5�]�a0�^y��7��"��|Ǐ5��� K����3%(!:�+�׻�2���>�dpe �ˇs�P�{8�⿾��'�߸j;T�#���Xw�
<���QE�Jߥ�/k�(F����`�i�X5�l}��}>�Áƭ�8RBq���'��g?Ѡ`���~C�MS��#��!�������+;�RUC�)��7�%*<��K���jY��mؼ]�I ݮ���9d�k�����J�(�iG�P\e��!�lт��/O&k	��b�$;T��'%�W���Ƈ)�;.X0�]?ߙҒ)E�ʡۇ�ms�d����x#ϙ5
������5�����jγ�.�T#�y?�{|(+xr���;��)���ϙ��S�"ESB"��׷c%^�t�6W�����_R $��l��LfV��1�(�&`�'0Ѯ8��/�X�}2��p�e&f|���C+X?>�_[�\�e��:�K&oXڰR�؍y�����MU�N���>,�饣/䷠�l��Q����\�(r���	)P^#*n�,������c��#N����^�^���&7b�Gb��-�|e����z^��:^r�ٸ����<Q2�kT��#Ծ������� ��� c��V����ښN����G��YVU� � �Z����E���S�����*����d��ը���.9���ȗY��k uv���rr�����DM��-3��`�����\H�@�w0b%��2����@���Ir�%Z�_-'��#�U�wH��BB�{�[�����B��J6��}�����H�,�@Wj��	�}����V;�gBP����A̆�leoNs��IY�/�˿5"㇄�E�ˀ�����.�2��|�w��g�VgA�l��z�TޤT6�A���53#i�����hV�l�/h�h�!eĐmC�9W���l
��l�l�*��$R�/����5���1Bv�u���`����i3��mo��A+.]-pm��5\�y�0�v��2#�����Z�������;yLh��v�do���l�V���WW�k��U#�t�/e�"�üx98��o�o:�掹q$b��NUrm��)ȃ)4�&F�ʄ�2��&���x�� �	�G�M�8|Z�<r�e!m:��8���=*�q!Tu�D��צj��W���Y}��V/K�7�x���&F��U��0�����Xt�����1��D��>��$�&��r��ܛ���E��߃����X�+�C�b��0����q|��4%�7�II� U�^�k��Ϟ)�O��J׎nD�Z]X���Q���j����X�K�S���b���W�N�Z�D�$�y�\Ko�!�����������ݨܾn>�v3������(ӎ^�Ud���p���R$�ԛ�>�
��`�h�#����n�_j�Ӛ�3���G"����.C�a �ueX��k�����i0�h������X���J�I�`<��%�Ǭ�լ���DMxmn�z̕Y�ȮDl儠�n\Sx�':�d����/�� ��-�'�+�s��B��"�N�Q�o�Θ«6���R�ae�E��_��
���Ӯ�t/M���!�ּ�
�&Vh�,�-]m�Ap���7T�	�ȬIh�藔	�s�v.O+���R���[���aH����_x���e=dh�賩�0EC���㋢�٭��@N�#�ǴB�T�&����6V�jy���j������@Q��Y �!Gy3������~�V����a�%���V����~�w�-x\�Q~&a�|�S�g\7�t. �eY���9'��Jh�0���wd_�g�u�j��s�j�!m֥��Q/�1�c8ͳ��m>O���'������0ݠ�ۀ��+�t�6������"p}[�7R|����"�s�[�>�e)�E�О-tz��}RE�1���~g�"��%z�,��9��j�gM����uO�R?2�Mӿ��7y�|i�����gk��Y�j���nY�g�:��u����;yg�%����T���0L��1���)��v��`	��a�z�$�)�N<V�1�Μ UF��%lz�M�'Vó�ߏ���},���j���2���0)��(�A�s5T��Z>�"=��'^�G�Y��e���ϕ.B�8�L/���K�ñ��9�m&��Χ���}m�H�¬�)7��
	�MI/�nG��$|�������_PD��v
�d�!p���%oaW��ޒ�MP��R�Z+�m4ri���b!q���_�?�޿�s�;�����"��̝��W4�D	�PA�*�P�_ᬒ��Ea�ob~=�(U�u��_k,Vsw��܊t󹎻�Ԅo�CR��!u}:�����6�C-�Z��!b;����եq%�2e ^	J�[BR8d�.����F��Ma[Q�t������3<���4͜*��C� /'a�P�c٣@@h��=�p3$����m�Χ�Wj���"� ���5��{�~��O���֫L�Ly<�G���pb����;�=A�fE��"N�-���h���\�������)$�&!��w����OGp��`�T��ImS��U��-���t���|�ؔ�W^x&M��`�,>��E#}A<=���ub��]��\���rݟ݊b^g)ɏ_�B������b�T�ε1�D��v8�E��3�h	��I�R\�E���!O��h��T� ;��!U��A{6��������_%X���0����DN�Uz�Mh
��λłhA$;�t{�Ⱥ�J�0���Q��Ř[�%�ʮ�)ļZ.q��:SXT
"\_?��}��|��c��WFC{�$�# �&EK�1c3��J�L�tO�a�l)@{6��\t�D�n�f:�1�-���fC}�Uf�>i���kCh�D�'YM��0��+��rȻ��R�'��H�h=[����_�=)&)����Gǚ�&���y U?by�����jwy]\��j���{� �'9Ǩ'p�0�_����|����O�fS����:�A�Ggô��zwW�� ۃ�������+���M��|��]
��A?a�J@<���eb��cb[dG�� !W#>8q�[������
l+ ���qu�RU4]Z��n��c����R�!��p���Q�F�k�	��X$��4q���'��s���u7�A�m
��
1��P|��fGΠ�X�r��*kJ ��}y|4���I��~2m) ��7�C�T�8���谮�|o_�+"~x�΋�[	�rI�a}ԕQl*���sG�ė�����Ƒ�q�/T�?Y+�p�&�?��ጤh�G�uo0���U���q���O���?^(�iw��JH���:�&c�Շl_���7���p��R�q%5]�KY��KQ��IJտ����}dP�N��s�+� �J ��RQ_2_�Ƃ�wu�u��1/\*l�GR@g�1c�!7}0!M�m)�#��e�b��c��{g�[�*�V�ކl�ʩ�͜M�����}m��;z���V~oU�~�ȅ:����Z�v�m��KP���Z�F��œ�o����gZ�_L���T��&���D|J;��?��+�kF+�~���j��?�DC�.y̓�>&��x(�~���ݶ-��ڨp� ��3
5�-m	�ܣpT�*B��+s]��p� �d��4�K����,��x�H���%��v��,������ŝ6J>q��uxӚ1�'��sB�?6� ���k��)?��"��F<�2e���(m�!���aU<�������ks c+�.y�Ɂl&[����2r��}�8���LO����ԭ�UO��E;�O�V�m��#��Vǒ��JG_�W�UM�`VL��.�|N�����Z�l���J�đ�=�����A��/���6���o�w~���� J��X'�C�Ā������Q�;�.y+���O��	�RM6Z�E�cz.����D�X�h��:�a�r���r+�u���cڼ]�9Q�����~�=â���T���G����x��6i&���2��z��H)&�����*�vnd��,(���Z\�V�i@��s[sǊ�7���+�J�F��ag����;�O|L�\�<ź
 Y\6d��
��Ӝ!�V\��Շ3�?���]��=m��V��7ܹ2��
�W�U����d�.?�r���2e�l.z�q�l�[���$ce�%*��:�M�!U9����2X)���&ՌB\��~wb�������>�eJ۬���1���7��q&��̙�`����.D߿�4o�S(Vt'����I��!� �[��5~�p�b�-v3�R���\]�q�9�`���F>ۼطB�؁5=:�RQ�T=�i�U��[���b�@�+X�5/����჎_�q�]c�ZQ�)9����Ya��Eo/�4t��D�;k]P���z}�D�!�E:���L1vs�5��y�2&s �V�"��j0��;�e�s%�����
O�A����\F`�X5�"��O��q�o�յǆq0�\R�/��?㻇�h�ؓo���h� ��[0��m! �{�e����h�H���4� �aA3�;+ִJG-_2V�㡘����+7θ��(�Y��`�� �~*���� h;�s
�"}���sS�t�2�z<��\�B��%Vͻ[�f�uȜ�*���ݎ��2d@wnԿ)�;��ׁ��Y�S�� IO�~ȯ�ƍ��l)�
Occmn]Ͷ��r��������cs�a
���Wr@��E���u.V6��G�WL*2�oU[KD�ul�@Y�X� Ʌ� ᖢ�ŝ���-�o	u����-k�d�%��.����RK�	Ƽ'Up���N�0$ڇ����	�@���O���E��^���*�8e���9�JQOt�|�z��&��u"��QMR2�� 1���{��� ȩ!���E-o�����밋X�Ď��:��_�T+0�}���s+s��q���aT'���vrl�Aɚ�弨����H�)��KUŴ1_�T�n�9�缒��f	8��Y�ǜ50V)zq;Z��X� ]��fަaۏ ��CUjD�y!���G���81�W�;u�#�<|�7pM�20j9�h�m�#p�����?�+V�h��oz[�N7�-E�O[$����~;C��ɓ��y*�TC�i+x꣓d|��`8<X*mȈ���p&9�ς�l�G�W$�k�u�p?�^��:O�-b�0�q2�-v�Ol�VS.i��y$�4��!t�Dom����cy��6�Ą��@�HƸΏ��K6[Er���4�y��V]!ye�GsL��)�br��5u�H����|K��<���?g|o:��%��>��y�Iu��
�D��ȇ̹��P��M����ٸCj`��l�&O��8o���O}O�}��:LZeC�E3����0�]��y��1�3�R�]>���
fm�ח�K	�PP����k[�M&��Wy��ù��x	i!�i���'����v��0��u\�ݺ�oG����բ�-̺ҡt�bD�T���T�U����#��V�,P��ب�K���;K�D�"�%��t�S6a<BH�(y�'2�됍m(�*�3�c�2~�	��|:����
������ ���bM���?De�U	z��u�B���LU)yDR�gIN� ,�n���@���Y�;��I}o��4����L����ay��ܥ
�w�]������F��m�s���"D�5��E^gmss��$�Ω�=<iލ*l'-������H��W�s`��S_/��&~��MNnD��\O�r�p{��ȐW�{�R��$P��s&/��i>��sμ�}G�n�8�EA'�nK���2|��1ꯠ��~�fJM�l��k����^$�f=[C�W�Ը�(:^��>X~�q8�D�Ϊ^�j�q�zǣ�UՕ�`�e���=-Z��D�-�Z�A���
������V�^т���1?cM��S��@����W�e���7���"i��wG����,p�xQNj�I�y6Ԧ!dW>��TN5��B��=L�M����T].
�N�%���
�x.4���h�X��Zupˮ��6���gg8.f��w�
���Cxټ������	պJ��ܪ�>�b��jZ`���R�Q;s��b+��"����*N�a��
�8z�SZʖ;���ƣV-�n�
�ƤHC�� '�"�gӗ©�Ptk�C��v
b�p>?�$�Tյ��s������k8d��E8abSY�g���X��)	)�[�ȣ(t�-&���l9��'�� �Ai�,d��ݧ=�����t���1���tD��9X*�FV�J���6UB�D�fBym�U�0>\m�B��ᙩ�b1vc���կ4I䋕b9�W��uD�,��k��Ћǂ8��`Eqv�;r�|��S��/�4��S��{�6*>������X!9�s��<��R!(:����/�����xC������'��MZ^��Ѣ�����ٹ�h� �D&᝭���綸藦�5$�^�^N��⤃���m�l��ш��hBw��E���7�_/1�=��Z�ŕ��Y&�&��Dm�g�͑�RqV$s
�'�k%��J-�� #G5��XS�WU�ʚz--���w�!5?�8�7pn�eb��o���&f�7��;_T�%����J�i���uQ�M�V��m��`n�����H�'����x��o�ex��E�
E�d]C��2Fxm�O�W�0�=�(���3�� �}|Q̊�H��{��S�E�7�@ J-�tW��݆&���ɔt�*�LG=��o����4c�-��j�I<)�5Q?̬�{*�W�4U"�t:Ft�-pg�QaEZ��CK�}o�V�	*G��@e�%t��Ƙr��_��>��Ǵx�:��W�+j&)��פv]�}����.g���6����q������*�������Ս� >b�99�BD vs��p8R�R}�<��R�@�sM��L.]t<R��m!ק(��� �drii3���B.��22>����y�`�l�NO�.�w<@=$S:��k~:���R�I�LGI�窧���Y7�*����V�~���OjD�����-=9T���%Y���&���&Z�Yy�߂oë��{�cHi������z�X�.K$ƙe~�-�Y"���]�|SC��F#pCD��f���s.��W�.��ƽҕe~�ئ	��8K��9Mx�.a�DCR��6�w���!�^!�w�:l5������UxX`��+m������U #�&��Va��KU4ï������a_7hF+*�vܗ/��� ,�*�\7�P�;Ȼ���Z��c>�f�W�S��r˨���6II�9x�?ٗթ���ġ�a�&���X;����RgҫCS�]nbȞ�z��YEԼ3�m?��-��O׻�m��6�%#�~���S�iu�ϱ�9�wA	.���V�zn�ĸ=�Q�_H������v����qY�2�L��M��u��B��k&���F*"!�6ͣW�;���)qя68PQ2��W��D�7ݱ���j}Bg���/uX�%�p��+I*Y��^�Sy�
6֓U��fgB�?Ԕ#s�ʹ][�//UX/^?��%�_�y�i��9暃���� \�b,���+�bx<��ʟ^�ȋ�h�M6��O�9��(�G�
���g�o^���N�p?�xi&����h��TC�
Qz�;�5���V�J��A���%8%ѭ�%w��L�ӂ߇�ȹ��3��4�H��f��3��Iu:nꆸ��ծm¦F0?Y�m-D���ʱL�}�:q��ˇ��Ѭ��S�h+�~�86Б�73�"�B(�V�ߌ��R�8�S5`�w����ZN��r�Nb�[��t��1��s�
ݕ��)�t^g��w��C(���c�hW�Y8���@�ӕ�9boi�z�肒ī�gl���bv<���ް�&����T��?��i҈<��א����\��R�ԯ��lj�#��N�� c!բ�d��P�S�_�P�(�|���4��������-�(�3]PRN��<^ټ��6u��5G@頚��������y'��G!N�g1%,�\��4r9��ޮ�G��=oL.v��lp���R�s-��1+%,ǐq��#	����ș���9�w�	���G���s��;�,����f�𷃮D0�X�����^���!�?LK�k�F�QI��p���=X�NC����k6�X�
n�����	gU��J�2��p��H��hsx�W�AE�;-w���E�����l ٢* �Z���9l�ƭ�^2zĲEl9/^�ܷ��u1�}v�J#����'�/[:���v���1MV�����c`�,,нf��0��u[�����5����Q�c�J%m�#)�
���Y2�=����&hx������J(���j�vT��)�W�%�P�T��c�`m�4�kj��l�R�P�C�Y��Q^�O͇Ef|w�ϔP�%{�n��2�`ݮ4�5+i������g�×���� ���Z���m�T"6��å��.�9�R�H��ʵ��SX��aԘ�G���q�m�oXx>�˵l:������0
���S��΀*%��11�������� Ό&Vl������4��u'�s��������GY*{_t����|�r���4�,�ON�>�Sv�+���z�vמY���^��@�	D
4��m�%2�WlTc	7Q��h+<3�����TcMC���/�౒~B;�Ӎ�����W��@��I�an��r���8�ڇ����cP&�ʊ�nzt~P��nE%n�C�+ôiQA�d�R��ſ����S�	������5N8���i��b��S[�\#���3��J��ƭ��R�g��$�r⌾8g��1F�{�l����
T �g�g���PW�(9����PQ	����>S�����|ԡ��.M%��8��Oۇ���GT�_Mݫ�%-�B���4�L��o�R�pv��<m��D^\m���Y��n�I
��rI��F��)Ti��5�i������V��R�'F���	i����C�ݔ��xe���\�N8�Y	��@������Ry� RD'��d��e�X��\>�pR9Z����Qfi��*��ۡJso��x�H��8|D�Mv`��g@.�j.n��I�H�殚m�}pv7��K5h�%6j@E���d�u(t3Ŷ�qM%c��ۏB�N���o���1�JK�E�̤b�$+.^�=ɚ����@���q�	����g�%��$f�_J��1����K�&��@��x۳���P��h;g0����t#/�([5�<��8h��0�m�kb��N�zy%%>
�Ua]4݀�����QD�R:���6��M��2Zۭ���r-*q�O�`�e�"9&M �i]}�;n�%���1�}�U�#��7v���M�mUX��X\ѝ�=�)S^xW������b�e����+!	H�5R��D_�-��]��Y��k��P_d�X�f*6�/J�`�N���}��6+��8/c���ԧ�UZ=\&^�@�����;4��qq�TM��R�?XHpgl���� H��O�b���ڷc�%D���.��gcw��Eo�+����j�G��b*k	 p�饷O��#�>d�f|�^(u�w\�\"�\��v0�J ,J���c�O8�$�2�\K��c�w�B���G�z��* %'%B�b��{CsιSB�ƥa~Z�����EnyU���rz�PV��_�GI�~:s`�@͸?%7�R�f��P���`�wÌ�8�TdtF;'6�y¦D�؃��f�O�.1ڗ��0;&?;�h�C7#W�6%��H�x�	���o��*<����`S����4��B�|&f(�{������ּ�/@�dkb�D�0�E{nKG�D-����^�v���i�3��k�q����|M�q�5Y,G�#�߯����`�A�Xù�^v:���t|��Q�ºv�d�s�1'��< D>������AwHC70���^�EO�9���G1����Q���Fq�x"��z8>�mԡ湭^ ��G�W1?t���������B0M$+�R�^F�f�� _ۼ�	��F`���fd�����a��Z';���R��}~<�����#=�s2��}�O��������'����M����Z�y�&@f���ۥ`��[b��}Q�����G�7�0�r��ǑrI�E~�S���c�z��XŖ��& �����|9)�寇N�<c�x.1Irv8����C��^H9"�_#I����!�5~0�W��T|�m=w�>�`�@��W�|���ω~�Ft*���4����I���`���l%�2RD��t��u����[��]�T� r$T!�x��LT� �@A/J� #�?��;�\Ԩ�п���,ם�^Wm�"��|�3Me����Rx��N�PǆS_���<;�'����l
>��H��0
$1��u��q�������3�`D�{ lu:�w���c,!���I��nN�䙷z�H�����:$�(�=��\��IB-����t�Q'R�|�+�����}��d�?�Zf�V�ˇ�ef`٬&�)���_|� U�z����9�L����yܘ���q)��	�)�	��m3����;B�5-�$�w��o���}�$5�ٹa��x�gn�!��H{x���(\ G���Eu���i����\�]2A.ݺ��q�5��c�ܪ��&O���<��_��X퍱&�<RK� S�Q��.[̒�J_ނ{�l;А\B�G�7�,Z�WuqQ�1��L�ez���iYm�Z�&o��km��&���a�R�U���m�r�ϑa&n�)����z�_|�e�L��;� rh�����*���2N�oc�!d�$�:/?4A�aU<2�C�d�Ձ$ڝ1�)��C������?V7Q���Ʋ�� QPjchCj� .Iu���}�������3�gC�9��Ր�w�N�_F�A�E�,Z6yb���?��O���np93
���~��^��{_ ��ݬ�p��pۢ�گ��yp����Fa�n�&�ަK���r�j2vi��$H�i֊��=�T䤦G��tYZ�2�5iv�?�g�t�^��Hg�l5�9�����k�	�R��e�2�,�v�ѧ������b��V����*߄��z���&U
�sFcؽ6g�+H-�|�}GW����%n���y.`(��!�%Z��4z߻d�"��2��z �j��)����Z��U�����=��C+9NZ�$W���q�齖1�3."p)6��M��:^~�����TmB�E��?<�Ɍu��u�l$�E��6l�;�L�b�m��^Q��ƛ1�o���*#N����R�A�i~���Hݏ2&�[�й�0��?�X4齡�K����x'��,��ol��G�c��e���U7rΝ����_!j�~X��o��jBg����:%����h/o��l"?C}��j@�V���-˒Y���j��d�V}��6���A�eP��kӨkU[�CD4}�K�����ղBh�u��܈T�c�P�K�S�3 �r׸0�T��%OC���r� ����5~�}�'�N�n�.�(��W���Ԝx�a�:��	���Jr�m��h$L�S��IS�KN��L|���xj�A�Z�T��Rz��e�U��C��Tow[�,��kE�b��MIG�]��z���	t���H����5��훥�_B6Fkf��v4D��V���q8o&|��3��;�(39���ѝ�M��y���"	��!��헷`_.E���
�e��
.�U;�/3�l�.�Υ��2���c�{W��;�:�oXSG�M�!#���Z9;���_X�h�,�|�� �n�X�<P���W�}%���b��$:�*�'Ng�V�@�Ϻ�����g�+�h[�EQ��M�w��z�L�H�����P�D�(����?��\�5Iy,��G��ڌ<�Z ��Bc�*�؄a� C
���M zB���)��Je�\�j�"��K�{;E
�,k�lKX#,٫�@���jN*��HW���΅7_WjyL���)�
yB�8�h}..v۞'[��M�Wf(�H�|����	��2���Y��Ar���㵖�y���K���4IQ���/�NP��<}�n�Tۘ��^�M� �o/��~ϜE\�;18*�+:�OY ��9��^���:S��)k�� ��i0�3 >6j�/�x�Oj
[8�YD��}�%�37���!�)3F��
�5�G(�|S��r����!!��"�݃�g��Z-��r�+��,�ժ��FmV}A���[C�P~��|���<�3X"��nw�<\@�j&5<��'n�����a��~���jɥ�і-�m�v�,=P��j!����Q�o�]z�XT�7�{4^�����V�`����/��4C�>l������\+�$����`�
6g�C�}�TN��n�;i�_����N>��6|����@7�!$��T\3�upz)�Bb�� �k\���ڻ��0�=V�hD�3��M��J�q�����ST�����[��i�H��������a���?��8(�Z~��L�yͼa�ë����
�7y�&���n(3�\�"�#�VÜ���پH��Y�� Y�4E���v�]�?���u�==�xL ���>���#��((
XD��Ꙝ>���PrmAt�`(�6�r���������=�o�Ė�.ߜ����d��d��w4ơ�z-��P|���Հ0��³3@1��@ �϶$=L-�0�mU5�G�S�J%k�+�.(�f�V���2C)B��fQ��^�����~P��Ѣ�%���)��a�üIX�N7��� 5�ց�@\�����85�� 9�"�d�	�a�W/�"��:8S
��|Bp�� n������3��C�e�p���z�^�Б@�[��2"��1��-M߸B��]�+_�l��O].af�M�95��Ƚ$�g8��4�\�[�t�@�&mh5|���$5E�x�%�R�^�М�N�K�J}�Zj���� Z�
!I���2bm�/�p���{�B��ޭ$-�']�$��X�̼5A�����dt��>�V�(��qQ�t ���k�?Do֢a<��8x}��ܚy����ݒͺmչ����1���!񡺉7�:~��F�9#���<�v�m�t�-ĻՅ�eB�ꚵ�r\�@�(g'b6����w�O�Q<�`���c'�e�x��b���X�N���vZ��?���s��)оhm4 &�Ͳ��hi
�;�5E���7�ϴ��р���1d�<Cn)�o�dwb+��=�?1�꟡~�2�^+����'�sOM{-[�G�3~�E�ѿ�s��a�y�mz����[ym�
�������8v�`:�Sbhyx~���i~�t;N0�P�2-ȏ>��^솂�<y�i��Pԫh��]����+]G�u�bQ	`�z�P��UeVb� ::/��P��vґ���ƊA�0�Z$?�<6I�N���#�n�0_�e.{tˑ��RG�TW�73�HE�[ٶ�å���j_��1g���7p�S*NeĲ�¨	���h�^nt���x���� ����t�[�A���9��09���:�SBP��������/�$�y�p�YT�[�M{�j�"�%��r�6��zZF�߹,�oZe-�Y�$��6�N�A�7�\��Ճp	�K2��EK��b�#��������Z���d���c7����w�Y�⺶�w[��6��7��'H�
��-��4w���(�����Z�j�����Js�e�7��u���g�r!^��?6ڨ��Pg_�u*����O�g�LJ�|�U_T0Y���(cú�S�b=2ix�G�M�!�>P�����9�Da3¨�$i�C�y,�1���'ʱ�5�������w�iR�ѴJ�38)�ٛ& ^�^yL�+|�B�&�J�����!/7���T��wg�(�ġ�ݍ��ؓm����{�9�/��)��Pڎ.u��r�/.(g�m�l��l��Ԁ��?�<�X�!c���"�39d�Щ�F�рt,@��^(��N�.���ɭm��O�^:0��c�P��[<���].��ԣ��|(�94�8�cZ79�ɣBYa�7��́�XWwɻŅ,���8��0Y������e���2�,�aV��ъ�x5r�)��)�df>�,�Y.�q2�"�#�!��*'���t�0�`���}#jo����S����v�Y�a�(VH�8��u��)�!ҷ���!	��i�'MZ�j��,��γ� L��SH�O؅�R�����x�@4,{  r�T7S�U9���i�2���@Ys�%Yu�*�Z�����|S�n��%g�)�R<K#�&�Å��8�;&04��؟\�;T�l�Z��Jg��k������0�=O��r�5�����]vkiL��(�lXj��������I��X6�Y*݁@QD8�iM�Fwq�9~j���X��M1.�<z�)�~�,�,�MN���=)r�#�އa�h]���[�ڛ��A3�>�7{s���9��f-*����e�'�I�h���췍dF���j�0\`՛��f�q�mw��r��8��k�m{�j��y�\�o秲c�Nľڻ��1�*9���ϐ+ȏ�.m�^��૮��ңs�7�C�h��,���i���`<�w��yt��$�,�6LϹ�Ke�=(��ᐋ~9�����D�g�}~(���/1��/���x5�cu�R�_2���f�O�Wp�
�j"��P[���*�Bd�39� (Ө�ᑷ����������)��	e��Dvfs��ς3�L����E�be��9`�� v���5���_P�6�� 7����S��IuWo�
�* �����X�Lv������[5��1�m�z��>ͱW�H�e�W��yr�����Pj��Qvѳm�o�^d��q�f��^������\}��v��d'�����{Λ�dx}wLbС�1���S��^��� �og�ċ��1�bRC��އ����ι�V�rJ�%O���B�;�Rŋ�os� 0F�<�~ǔ��|�wo0h��Ĕ{�uni�!��'܅*Մ�܂7�r�N����wx�o3��	��k�A���}��;mBP��\�u|0g:�т��Z��;ۣ�Y� k�!-&��T����=���*�>J�΁��t����pN�R��ù0c�8�`J�_u�*6 �H	����Fj�pC�8�D�?^��ϑ�+y��0pB�	��$$�:H�E��bk�
?&6�7�*�[�-��jkG`|�R�k����kN���Ĺ/�fT2�	g�/��<b����9c����RY����U4��eh�C'�O��M%�xDߚi��Vg�=���13���s�V���t��y�=u�o�~]qv����V4�8�r�rm��wx��4V��hH�X���r��ۏ�C���1�&j!n�����	��/���~�Nߜ���R<#Qj �^�#>2�'�W�0���u�q!�F9�HW�z�x^�+h껏�F��`�=�ZN�1��$�����ފk��� �N�K��#s�ܨ�^p�D�3�m����5�
�$d��i�����������pÙ�!���g�d�T����V��zY14DQEMvϑ��T�����:+9�U+���^ʒP�t�����?޻%��1�+� �h���FVfέ�l����@j��f�B!��5�ߥdfˑ��_eV����K��U���c k�3�
W[X��7d�Ow�MU���,Y:�cB���X����1�BY]<���v
h�a�I��Ie}��hh,�P*p���m4"X���3d'G�8g�6��6�c�~gx�X��0���LL�ȓ��Ҙ[��y��y��#}6��5-�b	�Cg�O�@�DM�+
�!	�s�WT�����α��2�M7�����3!#�	"�h�A��#F����~�rlR5�H��C�[�K6�{���2��v�o���f�����k`�nW�/D��8�-��K֞,�kB���q�`u]mg~��C�DT��{��g�K�Û�=/M��O��o�ܟ~�K8���n�y��њ��]����/M3��������H�YG/A���[�������$�O��\e�́�JcvN�j����ӧ�Ϻ�s����s��,�] ��I��<����aUZ�2�`���k��݉��x8�) U��~gC�]�(X=PpQ餦�Qп���.�����av�����-���ξ>�4~�H6���L��g�m�c3k���I5؂�V��u���C��97����z�h�K�S�#�ފ�J6���u$�T-�DC��ͱ�`���m�`��h�<nV6Y�V�v_L�N����I�����h�D.L.��I�v�K��é�E&����NwN��?��m�j��^�f\3̔��}�ao���]�<���W�[�o��Hd�*Ge5��^V��V�}.�VM��~�{8�)ãψ��:�96$ֱm�rb�Ӓi��n����ñ�|�!���jy��^��nW���:ɺ&6�~Xt��q g��xx|
V�~���?.�.��󞁷�Ɛm�ַ\:�qҕxݵ.'L:�J;^��g'�����[�O��=@�_����uu� ^E�s������'�H��ȓMl����)P'��8{g�u8tNz'x��K��{��=�Hbr���>F��dE���r�x.�e=�j-��e���ɂ��S��s~����>�����6�ʡ��d�斚�Q�bԱ:��m�����_iG�@sI����Hе����32�rB�&����G_�._�1��[�� %�W|�sŮ�@�е��m!�a��cNF	��@�T��t�N��4��t������W]��{�G\�c��"WU8��������� ys� \X���u�oȒ�!���a�Ё\�c�c��~�v������iʭ��a��8t�$�Xɋ��M9iFKBF�2�d�</�s}t$��M��m�]��Ue6}}��	��d&!��R1�F�pO�3
���ۿB%����rBֳ�;�q�ui�Pi��;��aϯ��!દ&]r�$G��A����#r�Б`�8�U\f^ȟ�҆]l��mP��.�~�z�Am��#Į$�M�LCe���ur�'�o4Q8���<��uv��eC@X�;��D+􈃍���P�1_sȰ�)�gXj:7�*ܷ��SQw�H��K|��U�h�羮1g�S�_JT��k];_�f�~�V91��u_;2�iP�N�-�$# X�~�Qv�:鈍�����f�9��H������Y3b|��2�"��g��A�:��S��xu��8��U�`�;���˨u��ch�)	f���*`͕y������ѸY�T7TLC�P;��`��%��M�Af�Re�A)ۮ!�����.͕�(e�3&�R-k����Xd���wt&�T��.w�t�Q>]�`������y��"(��l<+�y'����)�䳝��K������O�Ì�;8'\���ve���V��e�z�a�I����'��e���rc��9�P���g�Ȏ:|`"m�#�;��;+< �>�)���:���F��*%�^�m@�r�J�Z/�0=���F�<�L�w�G�m���ԥ�͛�>c��˙ؙ, �o��_���������Ҭ�T��l%yN����zdK���Q�����UIˆo�L���_���^���^�����hŵ�~O`T�I��� W��nV$ŵ�J��r��g�<�Ф�m�A#��&�i�i#l���[�z�B�#9�߁J��ji��9�A2ʲ�yF�2�"3W�K��r���+�\TN�Q�{�����0�gj=���!���ϥBA��b��7e��}�D�����^�@Z�+&��?�(���7qBĨ�*s��W&+���}$�0�Ԙ�w~V�MX��٥Yq�u��.��:B)�m��� |���l>O���ۂCG�00�R�����@���_!�i�E�߳��ש�5�-͈�.>2ɣ$f1� tF8J�ٛ�p��F꬗I�G��s��[)���k�|mW]�D[�J1˜��ek`ay�G����cڡ}����>���%TߥAg�C邈�t���_i�,��Q�<0d����	E�5��n��61OV�������p��/�Z;�/����+{�m­������/��m�[��.�N\ ���
85M�y[⒈���~��9O�'#�"��-�bx����5�9�n�)��B�J�Cm��e~�}M���M+X���F=����0k1⵰�j�4�_�G���5�\�I��!�:Q�����M~}N ��i��B���u��@E#a�}<EH� D�K��[����	�V`M(�oM�D>NB��tR��$䟱��cf�/=���]�~.��Y�M�ŦD`Lʓ�!��=X>��HW�!��j�sN% �qM"�SF?~v}+�h�ǣ/YJ����H��n�btyZA*��w���p�m�۝�ܙM�|4R#i��Ns>Z����<v�O�a��l�M�II�Fb�єqw���9 �S��C�@?@:�P�NIU�$��#����B2<�N�O��M��K�F�}
{ߜJ�����f�X��OoG���nyb�DN'sǾjᑻ]�3x6�+�����n!�ZS�c�η��"z��!s�RaP�5K
�����/*i�7C���W'H�YH�y��D򕯳��|�o2�<
���Q\ B��g��c��Y�p�{�&W����ʑn�(_�E�����%r�n�4tY�s�w��ͩOK��?v��S�Ξ.�����&Y�:	����i�t\�Q��i��R�CƟ$,sY��ӺD����&�Z���{ڲp;�KҔ���(��o�2�����
l}�C��}mC��n4+�����������s1���傸:�l�x�͈I�
���c���ҍ�e��=����f���(�>:��% @�OI�A���T���PÊ&��baj��ݞ�檲�[��&�^�O`��|�k�L<9��"�8.W��a�Wѐi�k{�1,fs��c����9 �t,����A�9"�[��<�+��w �
�/��aRR�wM%Q���v��b���}´1BuF6b���g<y\xi��3̻�a�L�

�g��r,�b�mi������t�!�h��5_��o�異����e�0%��em��TZp���d��l�����r�p�6M�j�>[�;H�w.�V�ʻo�%�\�/��p(�*�*����?�8��(���w���=�H�����N*�a��-�w����)T򮰡�]��y��:�����y#OW!�� ��ŭk�8>�uK煭e�!x������פ�@
bY��K���H�	PN��7��k<��b��h��M���i	P:�}˒�7vU�7��������C��'0>��M�<}��U葃��)�LQZ2��EK��������VN8�dp�3����xU'ئ�&kb��zΘ:��T�g|Wh�׏$�g�`d:@�6TnE�taq��"D���&b��b��S��L��#0��Q��8Km�Pm]�$��!�d!0@�K$T}��l@�1�Eޮ�Ȉ�f��x��a�tFhv��n41m(���{����9�:u{���������aea�G�W&�]�ظ��2F��˨b`7�i���(�0���âP���< ǌu/�|Wx��0���q;�2Rc`�F��?l:HқOI�?�#�T���c����[�f�l��'�cӺ7J�C6��|���nW���;�|.�N��\l��Oޫ����Z����K2���<1�&��gŞ5@�:�-�D��K,���sI����-Em�H�E�k%Rk��o�}f?�ܮ #��1D�W��ګ�W��q��=��tչІ��)w��_�h��2���$D;$Py`Yg}�?�=�e�����4�K+x��Ƭ�-!�LI�40�N�,B3���.�i>anԖ��`rI�L�t�*dσ�s+rqj ��x�bA��*q
v"�{�$�2����8��o#r���\6'��c!�gy'"�ߝgC6}d�#\�M����{�����:4���qD6�,3$q�c&Dq�+V�Ut�X�ы��
$8���k�լ$y:�Y&���յ7���)�eGi[���k���RY�r/ߢC?��1�	�G�?��oY+��n�f��@7�kX+m����4�Q�Ycf����?ݘM�y����+d8����=wDϪ�5|_�qZ� l*n�jigU�7�R%�W��-A�Kd�hp��N���O�wwQ'�sW�3��<�u�E�p�=_g�n��*�W�_F"�s��:
W�
rq;�P��k�6�(��GZ�"�_K0��
t���������iƫ>&�?�6�(��X���<O�7Kf:�w�_��#��.#�F��9t��I��-�W��Vt?j���"�S����f��j�"�XH�韗�zP�!�ndR���}jVử�M�|�4��;*:�J��?����Z1y����+��Ŵ>aT�!Z�d���4���*�3W7G�!�^!kbM�ʹ��N[tgg2 �o�%��^��3S�Lh�P�;��`�|(ѿr��8����ђ3z��S|�v\���"xW�N�d�$�ȹ��p��iKհ�Ô/��~G5E�P�)�S�gT����#���3@�׭sW��J�oB�����P��nX�t��M-��O�h��3Q_r*E�<���$8}����[���wf�Ӆ���G���[��fKj
8>�����J�6�X>����,;I�>��br�B��ja�;#5�G��T�L'��~�İ1;M�ݖ�|�UW'�P��֪�[�������A j�e�A7�x���u�+uC�����1S[��|�a&)�_�dhrR�y�.ۥ���K-N1L��1�kˤ9��v��).8��<N�Ny�*ړ��=S*W�5�TQU��Eun�i�x��@& +��&aQIx���WH��� ���˷w�i���`8ZT�LvLR�{".��ǵ)3��VAI����U�Tf���6���<�R��`�5�OB:%�9���14���6�E�j6�����n�h�~hwg����wN@��-s�T�q �O�����5��`J�F�gh�:�46|ӟ{��6�Ѡ{�Vq��#x�H����z״Ȩ�e�E�{q(a�"	��\�j֤6�h�B�{���<:��	�xD��79��^�p ��1�+~�����F�)V�j'�?���<u�5D]W�-Mr:�<����8*^���	�*-:hA�io��N;@��鹝F���9��ܠ^]��@�S-��s:-��?�#i󣣨EqQ(����E�)q$��}t��gur�8��=�*�-��eף��&)�P!=N��Y�p��C��W^
�X�}�`�]�
��^�(�9����w�U"����tD=�W1$�w��\�
p(c��m�ʙ� (ʐ	Y�?1ҕf�X쩍�"gލ����؈s%��ѾQ�8bO�zb����I5e]�������������bZꎘXV�x��3�˞�a����v�d}ƌ��%��1:�qZ�9�laAAp%�"��'m�!2^�zT՞��;��#�U`������Mt'�6�=˕�>�M���G(�t��;SD�L�S��A��ݚ]ƊsA9؃�f5<2e�,�����ɱ#�e���i�v�W��X�sbFS�[cٺ����y)�wj��g�rOM?����:Uy�P�=^U[��MA=�_��Cطn��z�sŜ����i��F�Q�_>=�k�*U�=YXA��|.̰/�k=�� 8�p�dG����#�+���#fQ�"-Y�ݟ'F�"�b(�(���3\t������	��*��oі��8�2Y=��-.@�^��3��q��c�X�
s���kK�5�Y<o�x�}?�#�9�Ub�6��9q��X[T�{à��~�YA[,�U�m�ܓ��dC.J�����=_�x9�gt���X^`�,�����u��6�Xy�M�.B���o���;kP
�%Ba?}��z�!8ZM?3�p�D��t��{I�f�bge)<��1���mZ�'u�پ)���շ�XaX�/,��(o����s��K�5 <�@-:�fw���&^b"�8�ކp�>��#@�-��}��qt[�ej�'*b>���+=^*pϲ�O��c�\���z�I�6������?v�}�<l��+���b=���-����Gc2�1�4ް��6��S$��ac�~XϦ���������y��n�ޓ�1!�&1ʁp�944�|����j/��K+LXXzY��n��,rb��I\e��G*�W�7g@~�l|��9J��k%���]�����0A�����cʋ�X��3��Ҝ7�dh�h�<�Hk��̞U�J���&����`�D*{j���v��h�,[ ��6�'A%$��8�4�+�����$cd���Ȭ������+�j�t�# �ۖ K��� ��x%��6�SqUx��0��s:�&��?�Y��]��o�'������~�麫i��$�R�eC��C�.� ���۾P�8z1��G�T>�T� &�Vl#�u4�_-Pc�Y��p��Z���c����#���F4q4n���Q�_?��_m+�In�3,��<�AF��e��s�L"2]$?X�"͂ў�Ut�^Q�dq!ƫ`W�TY����=țT�>�-�*\�/:�܎�2E�	��$h���pa
2F�%u�(kW�ϬK�S77�Z���2M�g����5�V�`�+�|�L���Z����f�_E�ۀ���!����?�z�m��B�� �VzwtG�����e�{��jcȴ�C����^vV@��
��K� }`�2H�Y��_"�լ��BW��,|Zc�Pw,s�%18N�a�j����=�1bEQ�
�Ii��7�K��%��(�1�A�ܶOo�槬��[o��emW��CS}PϾM&��ʝ>&�?����9����.�k[��ӣ<˻�`IJ��U�<_��}��*��;�Zu�Y�qLq����=�&Q�?��������j��z+�g���wݬ��d.8���C��^Gf^�9�O�)'��a.�1���T���J�L~�[�ز7���TXpʉeG�8�3�t�e}Dm<��i��S�"���#�+�ܛ��Z�W �5���OcC��C�s��xoO��U�I"�?}�� #���M�ɑ�۞ ��&��@�w���%�>�hB/L&�S��h-Y>�'L��yMp��%��"���
�&��>([�^��
��/��a��%���5�KT[��!�^01���������gaTS�2�%W�8�	*b�"�:L�w��zSe�ʹ\-���{�qVL:	}p�
<b�4��kL�.:�N~l�����2��D�Z!��s�9�j�篻���ٷ�zVU\�e���=E�� �<(+/V��g�퀩���%�ۤ$����$_�P�k<!Q����������2󀰛	���f<7HRA������"R㽟�1��>H�*�=�6���9y�q�њh��D�Ǻ��q�y���<ѝo�-�4>��Ka��:N�2;��@�P����5��0^�aa5�F�,)����Z��������z�a�1\�G�3�*���w���jv���KM]���+7�i�ʋWсIW*��1a�����B[������'s�~ڊ*z��#a�������bFJ�uҐA���1��ަ�¤���Vʑ��wO����Z1�h� ���V�?2��ķr��R�?7�ʿg@��[�O�r7��15-p�e��� �����������(��"�!��>7?K�Z���� �_zz	����-�-rQ��-"iz�KC{���cL�P
��Y��M?���9<�:�Kq�r�P6��4Bxd�.�e>Ek�C
.��y4�U;���l�Cz����1ѣ���`���~��z5,�F���ݭ���|-�N�4t~��ݔٻ`U�(?)~��WkZ#�	�w����i�ѕ�9�Ү��f�_��Um��y���5Vd�	i������9�,�"7�r�R&d�GoҺݧͤ����a��������'�X�%ۜY�[�@u�%��}�Z���9˪\:�T+P�6�O@n���ڢV���7����#�]���[_���F�OT�J�+��*�:ui0!;c`6Y���,BI���q|`C�;��C��$�ጨo�9:��ꨛ�{��q�E�T��(=��Kd��c)i����H1A9D�\g�v~�����
Bޒ�)�H|����0mJG�S/���6 }�ǻ���O��(e�Rw�^��n~b=G��0y��D��ϋt�  c�;�fV�9���d�߃Du�����Qwj��3�s(�`}|z9܍�cT����2"ܖ��\�Z��`#�bn��x�0�PӬ�m3q㨨�R��%�f�*9���;;�W��B�,���+i�����Ƈ�݋u�@\)������������I ���d��n���]��H�8���dkA�x hj���/3w���a��Z���Kɢ[�=��%}�N�m�����E���:�����uK1�Ƅ�!��WVa0&� ��mq�.�����1�����4���u鞧�P3�{5�b���t�h���\�.�t7>��]A*V�D���}K�eq���:B��6�;~��T�2bQ�B�Og�Hw���ȴ�:#F���s��<��Q�p� ����P����\<(�n�Ƥ"3p�)�4U��� �4PƗ�5��%�E{�綟��xc�j���W�F�L�3+N�F�jgK��A@m����^���^d�|b�i�VeQ�(�,Cԡ���B��r�UM:�V��W�4?��K�wN%�)b0�CZ��f��J]�;f�դ��m�ӌI�I=�i]�}'��W�~-��i'_�@��0����|V�BxU�Cz���~G��A�4E�l���Q�F�@�,��+{=��w?Z;J1${��q��+�bw�rF����A�ߧ�`����$!
(��l�ǒ� �Qu�߃�,����%_>�K��K���;+����"y�Z0��J5������S`?������Ņ_��:�z�� lK��:'�k���-s��$De\���l��ZqJŊ��)�]8�\�S-�
R#$t������ac�@�"��T1�bq��a�0'�v�0d��8��а䅦����%�
f�{铈�:oʶ��;��n���n+�˥��j�f�h���e��I<I`�K�1X��;C�$���C�b`zDE �[ Si�s"�{�b^��>5O�(��:�Zs�$nq���M ����,>�����0{�4����)SK16����5�{<��8�1�sVv �͡4/,��ڕ�6��C���N�x�C�������S�YD�����#�w邳�#�T��x!
��/=�ӱ�2[�I'Ѫ��Y\
��L�sÇ%��p5�"��<,@�:��y��Ğ�[�?b f�G&>�e}aA�f]�ftV�~&�_ջ#�(��o%8[ز��#p;�	o���'!	\88L'V�����;;0'#��������:r�R��k��\�EC��Ɯq�y4Z���O��F���R�p��_2/첏�������#����;�l��D[>R�W�7Cf�ۥ�}OW�!	�-�vT��[wk�k]r����*�*z?�����͐I��ER]�݁�w����D��:_ �@.�M��W��Zi8�j�������z&�"I�H��j }���+;�n��[#3Ĝ[r�n�͗���BC�, �U�Bơ{脞n��Մⷷ 0GHb?�g��N��� a���?kd��~�N��R	�zXĪ65��<���P�����AN��6�(���Wk�*�"��>Uy��"��ܓ����"�h��EEb��Ɇ�U��o�!�d2���z���7>�А��â�ܩkx���X�$�.b�P�P��R��I� -�xR���Q�X���5�Z3�xKw�tt"25��>>�?�gR�2xa�����Ҝ����E��tK^A�DW��:�I�{��>����v��cv���g�L�ywMܮ�82	�(�smފڗ���"������F��㈌�zW��h���8Hs37^F��06?{�Hg7⛀&�x��)$����
qft\���vg�6�+8�E�X xlib�)&�qNj�J�/�{��4w�;�TplogC��oa����滩�d>��:��8u�e���G�r^�K���5A��W����k=�2Iڳ�qr�ژ�����\myWN�n��f��i4E����`zH��
u�����rHz �3� ���u�LJf|�w���sK�� � �j�C{��M̄(Mo��<�\��OH;A������V��ts�B8qi��zr���^�C����MJz�r�Y�gw���S7��Ω���,3��Uus"h�|d]gN�:֠8d����2�F&�Z-l���s�U��x����3>I�S��(�%~<Nv��<�{����e7 �_���j.��_ʞ;��_ÖcS��8��0�� r�?��4�|�k�4�CTT��a��Mt��q��y���Q���}���Q�Ϟf���1�=�X4E�֫����U�	�r\:�k��)O�d{L�V�nL�V�zܷ6ĳ�4ҕ,?���>"�U�hQ�6�{9̂��<��AΜ�����[� r��7+�gY�!(4Do�u�Ux4��W�"�Ҵ/f�d֯�����l8e^\�.�+ٻMK�ᏺx	�5 ��a(=�{v�P�]W3CZN�`pV��.�V��sYA����_��6[�;�+�I�ja���&��f)��c$����j_+��I���7�&mM�R����PL/2�}�
�8�Q�?����@�+_��?�V��
����u���,��\L�uT�¶]]����g�F$��
��'>o>�ɖ(��=v�f,���S��W�|V��t�trd^�e5z�u�(�ݨo��?��oc���+#'��G��k���A挩�IrV��m򽆈?	x>`^�߳Ʒdi"�d�JlT�04����y���U�,}۰4��5����/�5�^g}IްI��x*�S�CP��
(b{���E�Yp�ٻw|v^��zO&�դτ���rh�,���+MطW��|Z(��9�6K1A�I�E�-�c�M����|�]�m!��` a���Ϧd�Z�F,#$A�6)�=o�ʻ�:Ӊ]�Ν�����
d&S�P�`�2U������=���
}�xkR�y���.��R_L�4:6Ě0
F�v�ˁ9?���eб��s$��������A�]���c�I�_T`�~&���ɔ+�cO�輱%����0� �+Τ0�i�^r'
8�ς�k�I8��"���g���A����]����-�ȵ4ϔ�(qkR锄��e틦�������a�����Z��-�Y$�P%Jaԥ	R�}eL��9Dj�݂ N�{��A"Q��Bo��+[�R(dZ+�r��w�C�挟Z�@]鎏[�@�t��g�p��gF��n�t2�#S��m��*�<�'��~o�� /N6u̅�^�����}�%*ͦ2� �gJ)J��H��oI��s&����x��g|�� ��R��&"D�6(��}�V��YP�2�?��W��x���7��#�f��>�����PQ�2xLS��I��>̤J�-p��ޙɍ�.�0i�&( �������w=������*�ӏ�WZ��0���I%ڂ��o��q��l�����#,����		�X�k�w�ʾX"���2���3�;�/O����g���fNU�y#	g������+�11˪O{+��ᇿ�c������WKq,�� �꟢���#{��=���S����M��]�	z(��RҤp�Gvx}%�����aI��1�����4,F�J��&�e���~fGt�ɼ�BoT�g/BS@�{��&�}�*
ЯQ�?����(��~�:�M2�w�V��k/��/���Ԙ�G�,�S�~���f��!��B�j5[���@0%���{�Қ����B�D@I�n�$�/ �k{#�
�Q�s����ޗ\|�4$t��X���W�EP�r�}_,��iE�f?��p{Z((�����>�-R�h2O�e�}Z��oQ��5��rڛēس�ʓ�V��-�Á�AJ z��a�]@�/T&���"6�b� sp��Z��]�(�e]�W}ŗ�9TED)1K�&ڑU!=����fk��5��,0G�smM*�X���N�z|ϧ�'����1tR3\���;���v��v�i���4D�N>�������n�[�%�ڰC�7�pL��{@5<��ru�g+�J�?6��	�h�8hD�z@|��rͥ�JC��]�I�(-��r:�GzS=��9����h��A:&��4y��>�V�zG���U�aS�"�v��<�+�q��	TT��	�F�At��-3��c�?���f�4~��`P�'���=�)k܏�aﶾI�X�ؓ���nq�륝�nj��W�,�擂R�~���J�0|�7��>��6�X�M#E�h���n��B�s'�S��Xz���L>�.*�P­�g��B"w� ���3=�*mN�g+'6��T5n��_��#�r�ͪ�6���k{,�O�qձ��^��>�����ye�d���,������݋^�q��[�h�����P7'��.!O����L�5rQ�8���a
��A\Y�Mڡ:_E�p|vtq�-�(y �1�6�$��F�
3|sr\ �x-��{�ק�H���/<�/e�w����zb�	[�_.�K����ll�d�E�����i�j�	��:'s]E~�\#RsHve}�]�?=��x����薠��:���� �Km�����^=V��jFCŁSU�a�����.Fnn��uH���mK��B:�D9Z��O���Ux��,Vh����l��0�.t+�n[�J֯P�{�PI�{\����Z�xb�(1��"� ��-z}6��؞�q�6{vsE�Қ���PM���hr� mҧm��N{D%��"p�g5~��E!7����B���Fo&9:��wW�=!C�l/��] -o�rdN�N$z-nyu�K��4��&�j/�8�����Jr�$y�&ZC!��w&<RO�{?H���<��૿��R���#o޻�v�}����ZEb���z����F��z}р
���-l#RU0����o�e��/Rc��J�1�	 �XRH3��ZF��pGgewB��D/�R�慠��^9�؎8G����#K�*
�S�K�K���
h��.i�$���~�E��D�@Nr�*���6�������~n�����ڀ;<z����B��^p�&��\g>7�m����*�����VY	���P�e�.�z ��E�����y�2�?1],���i��S82j~�џz�E���8��8S�) 3E�m�&h�K��|��<#�X�~�]j{/U@�C����$.8�3.fN�n�\�ɉ��aRf�K�vz<��� ��E��K�g��[��!*��8�ߺ��6��n@*;0��&3.��e�����ЗXL�E"�r~ �0��$J��u�K���,$��j��D�k������A�Ƀ�ُ���pp�"a�c���c��^*� o� �_X������1\K
na<�q�\�QJP�(b�Gzηq��X�G1���� �?�_1R�p��3iEH���@ǑTX��[����C�m��೗M$��Cx�7� ˘�>���E[F��a�S�G�	��W&��=���A�C!��@[
3�yǽ�g�����j��iz3�aH
�����h4+��h�g�;��s1��>�F�b��]��y��p:�#���mK�^�����b����\������?��LF��E�/3z�lQ��H�3y�._W Y��+R�{Ng�JQ���ϸ�	�{���M.$�� ՆQ��^�G�/�����z�X�*d����j��CH��s��}{*+����ߴe4}�)h�>Q���<�8EגY���eD$�� � ��n2ɇ6��G�@E��Lj-�����r�1�?3����U-tF����WlT+Z���ʞ�=C�F�2���-����yX���z�q�ugMu�ׇG�1��S��nS`��d&�ϝ�j�f�������Z�(�J��hp�����:6�U�0�Y�p6��*ѻN#9j�)t���+�����v~��:U�M]87�f㈦<��.n�����E�8y�M��F�\�vŤ;H���`��]����W�n+��e�=�&U+7dvlk�����|z�F��ڦlwT��O[��4چgw%��~&k%�Ĳ�7����U��5!J��W�����|Q�,,H�-�t��y����=~���>G^�-�xZ��0{F���~]w�5����\D�J�����J�e�>�.�X�_F@~�[M܂�F�,¾J����e,�@ ���X�B���EbM=Z�yl��t�n$��ˆ��Ȭ��Y��ˊ[�>�3g���3h�<��ʎ���?���| Ҡg
��m(���7A{�G(�0��:O4(��s ���1��c^>Z�!Aݫl��~4���~E�V�#G��xq��P� .�Qʥ4 �����o�p[�C3L��}��|�5ZT��oe���Շ�H�$1Qe�|�^��*_��w��R�F��.��@\#�	�V0>KT�Ge-�LN{@�eZ��S����W����|JoC:�1�V`/Z*�Pr�U�r�x~�N�̨�~��OD�Ag���+�����F��	�LW��Lu'�~�n6h������]�������3�A�.������Ez��R�&O�%���M�$)�#n�0?��Re���y�o�����F`� [�h�7Jw�z`q���������7����rn�E��\bh�Z�l�^PeIXPꨘ�^�q����F�N��i�ש����h����䌽kP�ߕ�.�����7���r��z{2�3L��:���+���w�M�&uUܡ"O'Q�(��?�ă�{� ©�Ns�a�B9�:�"��VNSYu�����$u�m��+�bqu�/�Ao��7���3	(h�i�^�Ox�M�r5��]v�r�	�pK���.�v��z'����T*0�r7��?�Y�p	��h��0Z<�J���X��9��J7�QI�mz��Ts����(x���ۤm���ճ��oS x=sc�o}q;����@�D������t��r�^'�����H�8p�l�FN�"D�d�u;�^&��
֊��M�Q��fg����a�U�H�1P�9#x|��Ψ.�xm7��5F�1��z����e������]��'��ŕ��P���O!��aM�T��z��Sfcy,qk_�;}���@�{҂�#Gh�H��w�����1t�7�/̳���|�p9�ف���
��y+旸�z����<�.�Ӗ�K7��|�츧[��O�/���(1s���S'�J_��|�]�G"Z1�o>R�`����!�(/7�O'��b��X���/c��>s�q�_��3��ʐf�DX��w<������p8�(EW5g�W�\'�;����} �2���WU3=.�I���ҝ�u3����TEb.�|��=��<VC4��iΓ'M�E���3n
�&����7�;mH�GڱA[�mͪx��Yd[71�{���Gז���&��IL�'�� 6Z�߷�Պ�G�±��}18����K~/Ew���!t�Q����.�t��qlq���Pʂڬ��*��'���/�1�xY>�_��ׇ���fġ�����$w���m��o$y;��g�;w�"A�~�(���Ғ�f4� �")�&݆�<�,������%l�Xpp�QV�M1k?�{�o��ϕ�զo���:�|�XŅ�"ˆ�����[;����A,^0Rq1�)�\��!��E�T�GAh='G��$�ǹF���<d�G�R���`Nފ�k�H�_!:<�u������?�y���mUxX�V�!��9�~��![���@���Y�r����Em���_4��̤ٝ��nm���S�4�\�H�l��.�l�/��$������.O{���r�O7�'�T/
^�[�zJa��Ö]˄p�eɛH�~^M -ƨM4�'�6L�3�ב�T�����\L��y@���`����m��|���c�Y���eDn�L��{��q�4K*"���W ʛ�3�L��[T�����zH��ӑX���l���n̯B��F�r�Y�Cx$�>I\x��yUy��[�w�$�]k��F?S14��:��6S�r��ũ/:W_4:�ՀE�4)N���9͉����ן�9V������ۋ��i�3oe�����A�qŹ�U!�m|i^�T���.���������� �����p�t��Ӯ�E�6��Ac��L���{�<��j�> ���i���u�A6��mC��s��6�Z��_.���*�l��Q��#΍s;n���ݺ�bL=���8�G����lNŉ5|��3Ӵ�c��� �e�� ]��kR��G��T��&��"M�Y�ɚ�r�K��I֪�jX��E�<�=��Y������ʊ�\PS��b�Ǿ�"�6�c&b+�"�S���ik��+_k�;b������&�9��	�$Ȫ�XU��+���*�I%΁�a����5����	��p�!_p��2$z\�711)�.@1YXz�?��.���oJS]}�6SYX5_r�:�ꊁj�U!�r�>�����uQ��W�C��)^%�d#I�$�ِ</#������f�-��tZ���A�J�'�Mg�I���O[�|���Y�c�L �S�e�R��;0+[g�|-�c�S���i���S�z�<��0���_ 8�&i�)ڜ�'�(cL��S54]%���$�]�8<Ci��4�H�P����	 �J�J�X���Y:����W�L�B���h�zRu�����L&��a������)K`x67�ם!�;��x" _��#��)7��$���ck�^��$��Ʀ%�_F����1�OTv�¯yB舅��q.M�ˈ��Ɯ��v+vI%⡍'!y���\�o����Q���Bu9�Hշ<�]�ٖHh�4�pه�+�'!����c�6��i
	����	���`�-<��^JAO�-f�ᾨ ˑ��M����wy���u�t?E1<WqgКb�[���ӡl�Y������++�V���z�sw�q�K<
��L���f�	��J���	�LOac< �/�*�\��I@f�S�׫ݡ�ipJBJ��<��{-�]�:����|Uv�uK�}�,f8Ă�(z��'Z����AL�u�E�l�?�Ǌ�	��Z<�򌝧!��	9�Cn��p� ��F]U����S(�Mh�s��n�	z�����q"�^~�+3�5^�K}||�����@x���!��]``z~�Qok]HF;嗓*�s���c5h9��F�b�Z�LA�n���1ܰpD�Xƍ2#')��D�$�G�1��|G�(:" �Ř�Ґ ��Gڑ�I���.e<��a�������Q��<r���;�w���oBE��z�k�T�M`�V?�}Fꀨ9�����o�R�m7bAyB$�$k�}��\�z��H�p���I1��Ji�[3��Do��s��s�3���S.�����+�"�Z��W&���熈*t�%.!f�nt8�*���;m�#@���;&L�P�}�T�\3�z��k�ǃi�S��`岢Q�cq����4��N��<�!��t�����ˇ8�e���K^,}L���U���Ys��G�^��3X��^t6�ex.G�c n5j��nlS
w�!��H�V�n�N���qu\�d�y�o�W_k
uT�j]*+����$�Pr���tj��j��^X�ƽ<�9���%����H���bi��Xk�4�A�����O�r�~�'wnz�4_�Xl��S$
�� 3q�)}���C���	4Y�ۏD0�M�I'��y�29����wV�ʯma]~ȮDME�����`��ڀf���=�g#3/N�#%^�}Akr睼@�	9Ug��� � � ߘ�Հ]��ۜ�v�B����Dؾ��[���P�'<��Y����� ���ٷ��W�*~�Ua�`wPIW���>9+��k�6��p�i
���ʘ�C9�� J{�v)��V��QŃGA�攳�2��I�t���7�L����`4����>�T����=�壗p���:��9b�*�Q�6<|�7nf��d>���IC�7�QCģ��dx�l���&�3T�����X���ʿ!h,��k��D?8[&��ǿjǑc)њ)�#�v��	:��W���asN�w{��T���$M�3�����#D��'���@�.?ֲ��9S����hd�#mj�i�Q�����1O��ߋ+N�mX��4���1��&6S��(�J~;s�b��,�-�葥��+]�ԣO�3V�l� @})mo�p#��\��S\k��[K�
������`�f735�������v�u�9�"x�B�v��z�BB �7}�B�q�4��8٧j/�ݭ������;�}�MM�[�t�%�3bf7���{�IY��+������,�D͕&�I��t����#U���f�N,h�Q�J��7�w!C�yX-�qH�%Ƞ�d �'�s����_�J&��)��0��3�1?9!��fXiI�s����Pz�=��
��&��j�dSF���xu���8�pk���%#��Ul�hQ�]�_���֯��¸J���Ί��9�Gw�{T:ܦ����1��m
��`	[F���@3�N�D/V"HD��Ԫ7���XH	���bQ��`��q���S|^�3�m� Y#%U��/� S�N�ܧ�C�����&`k�=���m*ܑW_'��::���*���֜��\�}Y2����Ó*!���/1_�b�	�i��~}��D�?p3I��S#u���QE����;q��N�
6����ʣ��?���@�T��z�R��ng�-	�=�a��[���7��W��r��{}�V�I.^`�@��fvU0���E��\tO�[a	*;LhWƇ�_Z��+!��ޙ�f�L��gh�U�6{���>�`M�KI=�͍#Q�P��Gk��͌�/X{�JF#�w����.V��w�U�=DW����j�ik�v�=�ɓѵ�_��_g��z���@ �]��<N�ܭ,f�[�� �[��@�o�y^�WM�h+K�=?p��<N��aRp��o�M�F��V�&�n�ȎE�����Ia�i��V��r<�R���R���Q���6.I?��o�{ݣx۞��N�n�4��/��#/�>k��!q`"�O"7GEq1O�IK��'? >¶�ip~�~PP�T�t�ݏ�m�Tu.�]�L%Y�V��,��P���5u��f�2�����抅��v;v��Z�>�DL��M�&����*�e�Z�گX�(7���ߙ�h�W��j�a��-w�u�¨ܬ��/�џ�:n��@h.�\9�aҰ�K^��JQ*7�*��L���~��;��<p�*aLDu��B��9�>������ �A~�^�vT�<��������(?3юgur=�6���D4u�X�ʟ4.��T;C��>����X�l���yG�^>�� l.���i+E9�=�x.�d��Bi[d�G��yL�������ʗ%��A���,���ze�Z�H ��@/�/�ٲ�j��!w�J��V�c�{_^^��o;KU�z��z����i�%�:�-�R�3Qy�Y����|fx����|��n�2�F�g�i�`��n3y�0�=��O`xj�)�	~5�~�A_d�M�!�.�O\�3Ϣ@z�~�;2����"f���qA��/^�u�����p95���->�R�}�ұ��dA׺
Ȗ08��A�[>�~�A��Cl�U鷥���q:D�x�L!�nx����F���Q��ۃ~o���ä�[d_��u"o1��ӏ�7�;�A�W���V^.g�:7��X+�?Q��8���^��5�`��ʪ?܇�O�Q3B<Άޓ�qw�#����l����M\мPDծ|Ri.}D37/D��˳�.�D�]�P�j�������<7�M�1>��ρ�2(��sI�m��$�#Ub��&�>�	�K���9u]3���i(JC8����Y$��#.�*$��CN��BZ��V�lb�ʼK�`m�y�m_[�T)�絋�˓4i��
86�,3��+(\.��+)��W_b�-�ۿ��;3�f\�0����I�Pn��s��ӓ	֓ѩ�W�M�r�c�Cҵ`����,��e
�8פ(E�jK{A��eQ�L#D�B%�(��>�t��^z����r�9ۅ�i��`m�
�|�����P��� ~zYԸOl��F+V��'忨��3��6��#|ys�fO��_R嗁>Oo�t�6_]b-\diYA���e�o*�) `��  B������]��o�1�UXL�p%恫0��i��<^�N�ci�.^D����j7Έ7�][�M��h�J:���ip� %k����XCn��"M����V,f��1Ҩ�ܩ���d�K�YㆨA��Ze���c��E�V�H}e��&�]��!,�V��ta
9UR��\���@8ՎΊ�[3�P[F0=:Ӈ\7bi1HH4���,ϳ}�>��ж����8��3�I-G�1��U���\����Gn'��c�Զ��І���;"2�\����\���������+�˩�� ����?zұ�?:���
��bG���@ �� X�h؛?e�M(%}�S�V��f;Uj��#O/�y� ��?*�ދF8���ʷ�n��������~��14G4��3����ND� O�%�>VR�9R;���<C~{��k���/0CU�&��EU8�<Ή�Ka#m�[��JՐ~?5tf�4����co��\��LM�����>u-��p'AZ�m�����!�����`bz��&��cr���<�������!\��4Gx�H��=n���K�&��
u�a ׫�< ������T������h�cQV�( ��z�F���܏~���������L.	Q	Z������90,B�1�`-��W��j��~��7�0(NM�6�\|۟�>9���sH�2"^��i\$rm`?1$Á����T��Ǳ'�c�("M������H�s�`%X��k���uX&�H5g*gZ"��y��ql��rj��M]��������P��U0��!:�'.�õm���8�C9"�`2k�����w��	)�1G.Ɋ�b���-��|��ΤK�xI�lt�6�%����8�O��u"Q�V@�_=jZE����Z��H���|�R�/�������٪ޭRb�8Hȅ�H�d�
r'Y�NW�7r��l5�C��𺅑�2�Ȅ��G,{�u����2�����^0��E����,��26�������I#-cqTP:uaԮ�� ��}nl��˽M����Uj��H��� -��y���l�� ��ع(���%6��h�$���b�'cZ��=w#�-y��t�����L�����5.�֣&�Sq��lή(�fz]M��*:�4m���S�(��	�J4�����kv��!�7�`d%1]���#�8��L�PH]LS{��L)������w�d!�2��7�w����_*M��wG�IA���83n�"M�b�5"�p���1��+i�K���'��x�H*�~0�H�{Ĳ���W��h?rN�k��׿8ֳ��_ĵ���VSު�)�XBɲ3���ō8rO�[�����Wy��)��>�y��F�����&x�l"�����a��m0UF$�Oq�{q*ۂ\��DӜb�D��s��*`�?����|X����A��9|��?I�e�i��i��!{�����Ŵ���㫅��'���_�R���̬k<��{�-t������Of>���R����e˧XR=�5���y���Io�j�&�I��4b�����`��Y4�5��b�G�� `Q��TyO��R�k��6�ϯ��	f���`=�Gf��<>�Q,����&ZE��jӏ�l�gÑ6�K֯!���Ra#߬���i޶�`����[f��K����#��O�b#���蚯���%�d�p{I��2����H�۳�'_�Mvf�'i���M:�����b�K߫Ï:K�ϩ1bK圥��T�S6h/x.�z��V��.�`B+^���h�;��S&�8��1f�-�Q��,(I�9�ȅ)���0���.��Z������mn������X��|��m�D�WkP��ӑ�ٷ	�$��yj��~o3է�u��8㐟D�����^��{�f�d�=���J�S���dֶ(+#{|�D����2`ݵ�9���u����Q�D�9sq��l�P�n/��$��T�{�3*�k�R������Å��p�i�+t��)���JUEP'�f��ld���0!IS���s�k\k�Y�ב����EsHLZM������n�c�X���%�d�����`�� ��yJ.P�Up�`�Y���B�d�|zFj)���`��㫩��5Yfj��q��n���޽�e۾����u�e�´��-L�J\yeA����>��j��])��؝�Q�3�����	=-�ƸDC8���??q�簅��}����[ ��y����-+��Y�eC�������^R����8�g��(E:'|�,�&)��8Q�)E����3�M,���a��:����$�r<�O x�V��Զ�s̕9yq-$?��Y��_ ����9��|f9���!(Ǎ�UN������%v���t����bo����x󟚤���[EO�gA�i5����0!t"�ig��Uw �@Kx92�8;�s#1��������Ь�H1�F����?A�Q��S�D�]��@BP��)ؚi�sI��x����7�b����#�s�:T��I,�gL;HR�0TrZ٘��e����V=�w�.n�˯��'n����%������I�Ņ��o�c"ć��+��ǥ��j��wx$b�rU��M'����GQpl�j��+��ӗ�p�f}i�pҒkgk-6����j�<�n�m�2l���q�L�S%��GG���c�Z�6:�͖]-������_=����Ϊ/c��C�m��{LNF��(�3��T�<8��d����T�c�Fx��-i��Ҳ>@���`��t�S�GB4ڮS�j�P]���df29��QɹX����b\w��=a�" ��E [,_����> ���z�[C#�c>l�=��M����&ߙ���27���Q��
�0n�6j[[DMbA��S"�G�M���]m��_π�����0�ԃN|�I�����%��GW�։k_����� �J}�F��A3�9����^��ޯ��1���o�v���2C��Y��,�^�T%g�#^�[�(ɨi����H���+ɫ����P�5����!�ߍ�Қ��geX����`X�y�[�S�촂�Y��D�ֿOC�
(|4L��}�\L�<�	����e����}��3�f�R�,��G�}\���#\Oܢ�������3畜$d��)�z��NW�O���A������$#7�D	��,n#)��7���p�j�v�3F��K�`(F_��L,�L5Q��:���K�|���GP%i1�W�aw_�wÛ���p��ȁ��P�;p�L�$�Tu���gw�X\6���Ξl-)[�wm�U�D�A,�kw�po�����fH�G�������e s��CTR�g�xV�x]�T������ ����τ�;����jS?���O3Y�IJ趓Z�����z�kJo' ��([�/븒�l:���i��(`A��Me��E}i�0�?�?��:�J�<~�/�_�nR?�ƚś�\;+�$�[`�:@�`�����z�v�<���p�X�P2�2�76$�xGI��W�^D|��V�S򘀅�-�7S���^|w�꘠;���pt���/�ua�ÂL�r\��$u @ن6*��+�9�ܔ9#����Dp�w���4Ƿ&eq�)N[�Yi�̜X���=��<z���쒟̳���4+ې�����q���oG�O�/poܸ㑝�Y����ck�Ϊp����i��d��m�@܍�`uvp�	��=ե3�wU��d�IC�"��n�9S�hˁ7����ja$C-f�)�u���@J3Ms:Kv/#�򷒑'������ӸR�����\�lB�jr�t��T������8�c�����b�N8�������(͉����	�z��|��V�Z3c�j��Sd+#^8Q�{���<�|1*@���4�/TRa2�w���ii]M��K�Kr7���Ӝ��
���J��qӉ�s�tG:a�uR7���µ�gl>���vR>8��?�MQ�n��(�� _{����Z7|�!�Y�%+5�ؗrO�n+a�^l�Z�l.O�4NXm���;���<�������q�����@���DwFF�B�Q��Zw
O#T?����!iL�CaQڞMb��TA������i����|r<5�� 4�uH�Ǔ�`���3��oɒ����W�埦S Ι�����˶M��$��	n�E��!<�S �Z��W����v��!����mbm-0��HyL�b��W��lO�d>�x-�j�!��6�-�;>��T���l��r��Q�f-1�bd(��c�?	��{���ܛ��P��;�L�+#���q�ylDI��Pl�����d�:�Q[��롭�[��ᠴ�R�����@�剩
�N 4���ɚ��!�Uu��N��D�����aW���gnQ��i��D/TZ蓪B�?.�g���nd�^�Ȃ�0����B�_��[�/v�{����{�����v.��x/r��b�)�Mq����u�Y�|�9��.o�"�}��,vg���2'����+x�l�� �q��@��G"g�.�׾D�W������`��ׄ)�)xl��JL�\Vk��/�%�aB����  ^��Bز��q��=���Y�����_�7�U[�r�x��z�\� u��u�Y`*��a���N���l�lf�fg��1��X ӟ`Ț�&�4��r\:�"T���̤'3�[
v[|?r!Ck���k^+9V�3��:D�׎F�6��-� K����L��>\�Uڽ�X!�Z�$?�&j�붖�`8���pʵ��̵�f�R���x9�ÿ`��@2��C�Z�4�������,U�/�e�PC��FE:7�N��K4����(ފ�3�2O�hK1r ��}�Ac5�t�����O�3���O~���2���FIJVa�1���U�/9�t�3p6���"�=��_!拗�� ��җ_�wɆ��厱�����n�P�U�??6nSxu_����&�PE�Z�����&A�YO�zE ݠ����j`��o�@�_߁���Z$7����&̄sK}��bMW�|�;ް4;*։y��n�૕����w)��S��Fʤ�4��U�y��N�]��2oLt��/�Z=D��ώ�A.b��h�'��Q�%��9
;���x�%xtqJjHD�:���&��M�ph2�&I��n��fr-��±��MZ��!�)��8-��q^��V(����) �9|��X+�:^�~�Ug�a��!��U�&6�S���S@�,0�	'��iB����<IIG�4$1��lE�i\T)3��H��$P%כ�W�X����@j�l
A�p%9k{:Oq�,�r.�@��p]�w��oe`G��l��p�u�x�rX�P�x#�l
6�5��>��
���e���zz�U�{�3�$[��S��|��=�@���܉VP���ً�����J��Q����#�[M�T�LwT������[���qǭ��'xz~�0�[_X��^Qf(xܷc��/��E�~<�����$)c�4
3�o�h`��a�+�O*t���e�5�-����A[�b^��D� ��I�$������-}a;�?\ \�ѫ�7~Ƌ��BH# ܫ�Ǿ�7l�Kj�P���Aи����1�>�'HW<:�w�A���5�+0���RQMF�{���C&΀ ��	#-M�����E����I�| II�H�#�+��~���L�қ�9F����q�fi�e=?��cz��'VV��l(4���0s0��҉��ON���X�1�\�|�μ ����8�7��%=c�n����7� �z~�0�t��ȫ���%f��sκ>�KMO-�R�^�Xe�p&�MwBgP~4x���7x���9�ت:�~[����N���W���5�n~��Moll.Cn{�7��N>l/�}�Ӈɱ�v�>��^b��͔���tJ!O/x-���A������L���S���6�ϵ��s�M6�oYES�3-���嗽��W#���N�?�+;�t0xR�d�DG	ǀ́��(�#��S��z�
*SYBʄ2N�iokU���}�I^!G0Ftk��6��ߟrA��a�����ц�N�3)o����KK[�+�?����k�a6���� 6@���j[}�m4F�_�^4s�!nsK�y�B��;0��j�z�>�
.�����ٲ��PS-�p��y#oCy�\Q��<�&�O
�c�)� �R4O��7.��>�s��v>��]��P6V2.��ǡ�s(
O�Y���Ǖ�_">*�k��9�w�B�}Z��OkCY˅��'p;��{����lͭ�Gl����!���mW����U�З`�V]!���"sN}��':�(xd5'c�H��>q�R�g�i ���J-��MZ"h�f�AV��hb/��^�+g��k�UgEnU�)q�>1+����B�s���?"�p�J8R��2���ִ�O�":����'�Ck���������a'�/�dQ0a͊ >���7c:^?��M�Wm�k�J���ݯn.�3c�+��q�	r��]���N%��S���x�=^z	cy�M���P�Fd۾��)��ͪ{O[�Z�`�ؕ�Kc�YRI"�o�
W�')	��u���FYr9�+��=��-��X��x�a����ΟY�`�K���Рc�-�@�2̌�?5Ϲ����55�q@y�,��UA�LyY�*�,��r�]��c�b����V~�<��O���A f?�5ze�g@�ϺQ�%ɚHt�P����U���.4�O��r�#]rB^6U�N,�+����\�`C�1��L*���Ω�]j�+���~?�x��zCX�Ӭ��o�ĸ�9Du;�|B־L���i�J
3��}���Z�o�� ?g�����]z~�8��]>�L�r|��'CPJi쩣����s��s- �a�����E�P
.�9X��ig�+VL�Y�J /}P5�ټJi;`�JSk~p����㼧��l�*C�B���}ȝtrj��Jw�Kb�{�E<��:4S��Z��ED^?P@ͫ��7�; �o:\q�6Gw[�z�kÍD��$��He���>�7L�K<fFp�T05Pͤi�1N}OOT�@cp�xs����(�!0�g	�z-�������KLs�?5a�ӥL�)N�;����� ����h#�X0�P���Rb��L���� �zE��f_����XP����e���e�s�u'��Ƈț��Ё&�z��œk�{Hz�ktg�j��˂7�R,���뀐Ƀ�r�E'����!���)��b�U/ȍ@��A�~����U�D����¡��Bb�=\��5x����T�J�S �� ĥS��+����DDd)a(c�I$a����&�h�@��[)�/[R��<E{���r���]��"Y�x��2��0\��5S�b婇��z��Ħ?z�?(�d�[�,s�ݟte~�¯��T��{��vh)���f��;�8��{t�6�d��?CD$6�ZE�:��ʷϋ�5���8����Sg`X0X6̼����l7m�eO%�Qe`Y`��PD�rE�&�ePOj�\_�zfU��,�-�`p�8�����_J��G?�1hg*�����7�lXR�\7*��jT/]k�qs����1�Lֵ�d��o���I8�F%�dJʛ�o>~f���D'���ws�a�؏��<�d��r���^A�}v�^����U~֕>�ɥ�--��Q�NK�ޅ��UK�s��<��_�T9Z/�䉻��\���=T��J�m��b'7DޝԲ�뺈������Fm�2�o7��m��=)�� ?X(Ï���#��-�\�A��u�2���Y�][ú]��b��;�e�����}K�'VKwn$��7�'�%�P�GL���L<���2CE��n�V������L�����<d;_���r
l�3m|G	(r~�p^���ɍ��PϨ$��:/<ӝO��5s΁/ҽ��m�G<�`���Q�X�H��O�}��>Ģ�DIn=��nO��%���_���^��m�RW)��SZ�2Aoa��K�ŭ�7O+^�\�1ȕ�Þ��T�P"��$|��c0H��u�T�eiJx#8RAG)���/����5?��ӿG�!�ܱ�k0�<�:�+�� -�ݛ�%�MD�V��L��A�wN�+/�q������;KXhu��ŏDtE�����`�Wj&UQ�pJ|�C^O��h��R�1��G���$5������Vk1`��]ǁ�1�$^8wU��ݭO����E�䖝1��D�H�c��9�Q$�����3����p�a�{�geWJh�weQ�霧���'�*���<�]IM�R����;XyX1mm#5�T1�����=u���h�aS�%��%���&�#tX�о:+3�Ff��>*�ȍ��a0[�|��R<�X��a�1=#x�-�.n�M�p��z��6��S"՟m��0t{|��Ěآ����.?J�G�Jn\����$&�#�\r����f	�a����+c嵀�����p����~����kF�[�f'���1�	��]�����%������[��a)�x1z�m��R ӮZf�P
&/n8Y���#�#�4677�����Ӣv�ͧ�frޞᴍ`�
ó�RNKڷb��?�	A���MUw���:(�/�sg��>�|��ˡ��12~��G�Զ�M���a����QO�%���/���a�p�!�?F��r��b��A:����m�;�"T�ύ��=�K\��6q�r�ՈJ>�&���yDh��_�D��*��I���\Ϣi�J��`ē!^�F|��#hI�"���2^T��J�ԣTno��'OT��0	6�
"-�$	�t�,���*��1V�h�rz��jY�������0�7pG�3,+�!�o�Y��e1��R����]f�2��bH���	��BL��\�����=��=zY5S����=-�BC{ ���ح��ѷu��n��� &*�TSMSf�Z���R_|��c���ٱF�+��m�c�h�E
p�IaK�?7�W��24�+�� >�{IyD�:�]�C]Nzڞ�UfI'��� ��Ź��J�����O�qSy_��{�1�gH��uLppw1<��Ì�^�m ����S�}�I��1e�rM�MPW �r�E���C��{u�4z�8����$y�'\��| ٳ�SP����A{yX�A޶��bQ�s]^��f�����S뭸,M��G�����Ε]
Q.�n.��P7}>
R5 �+�1�=�l^5�Wrx�,ՙr{!��4/���"�sEd�� )A�`G>�n��U�[m�����$�<���N����_�ٮ�a�-��r�R��ViQ�N�{6)�A�Q�r].}bl�y��mt�/2᫟Gȿ���`ų����|�?��uQ�)u�I���1g [d�U�i�����������^���=&;��mC�\������Wx��fu��+� �T�}�#sh1���rކ���?=�k�s�Gh��I�-@,�~���2/b�������_�e� ����n���:��+�y}te��x�����
7pU�A���F	�+��}>���PRsҁ�X��#)�G��s�<��B"'Es����Z�m��H��ۃ'U���U�@�UՍX��G��(�bFK�8�����6llǌ�I���?W��\0%|���%�o�:-��pVZ��[`���c�.�� T��9�gahצ���U�rY��b���F�,S����ڦ��Tg�W�����" Ī����F��?����1� �d9_��%�^��>q�H1��l>(�Ŷ&����Ӭqu%��<�s��n������/-�BQ6~2�Fg������)z({毦q�yo&�UY�1&��c�a�ҌY�A~���?|�ۋL	��H�d~(j��tLo���5���
�8�����w�u��Ž<dz���_�"����0d�J����/�4<���њؓMW�bc���� k��ܭ�����wI�"�2�ąD��'�����<�=]>ӈ����n,捒2"�a<[h��������V.Նf�����j*�^����d��3/�+VPhjb[1&=5�>!L�z��=��t���?<�3��2�ԕ֜;%p~'�ɚ�i�����C�n�c(:1u~%4�Ud���%���p�yMM�ɍN,]Pzr���*�:��l�CNTJ����I����؊�O=Ƒl��Ѩ}6�W+R�:M���;�Ϋi�%��CX�l�8�;�O�l��.nf���$��
s�/s2")<�s
�D���Y)��e�Vכ9B-	�Ī���Գ`Ԝ+��S��[qFp��tTT	��>'3�\І��;E��oC�P�1�	h���+�V��,L>��q֙�X�^ŕag*�_nm5[���.�Cg���G�[<��-�4����3C��YMe7�����p#�����Jf���5T�Ɔ����(�Ľ(���R`�3�Odv�]I�{ROL�>�����/Ȫw���wꛓ�3mj*�oY�ϩ��3@�iƿ�"s�M���8��������o�N:�}�:��DobD�4ƺ���j��9	�1�i��2�fy�EmeÞ��h�S��|����A�M�k5�q��N��g�yѸX>AF��f�av��2���˂�ꁄ��"%�*8��\[�8����A���@��{��C�g %i�U��W�x���C�z�-/#6(��t5{�����]�*i%�G�����P
�Ŏ��vAy{�{��m�>��G璄�<�-�B2����l��N�3Hev�����6��JQK��b�.�63�ť"�hP�~.gު2'���.�v�}Ӷ�WI@R���w�I+�P����w.z�n��aR�w��/9��S�>&6���Ye��:l��񪈂1(�f���(_�q���_#���T� �4��3�nEw�1������ߏ$�v$`���]dS;zP�l��A_	�J�R��i�4�>����؆/xH��� �e��J����eB���Q���+9���t�1�5b�(XI��!����o���Wrq+�#������b��F�>!j� ���c"Q1��Lm3~���yUW.��.��!�L��v�L����)�/�hb�b�t�!��J`c������͛���V?�(�
�1�!$N�7�9oz^�]��9�Ag=%|xߧ~
����F8h?�9�Q����o��aW�X��:�Y!��N9ڧ�.>I�1	R��X%l-#V S\��k���i�Y`P'�E����:唝B�"��5�U���U��x�jц�����|��%?(�*�4�TQX8�M�u3:T�jܥ3�� h��D���g ��4rw"9S�.��&�u���:��@�ộ.�;����ࡈ�I^�E-�ߘZ:��,܌��	�����o��m���ۉdd���8a~<A��p�����3F�NK�5�BN/M#��96k��:��23j�,�2'"�W�1��d#�c:ܸ�h=�,I|��bë�7��yk�~�"���Pl��}����A�G.9���VU��E���� A���U�0�y3��&��w9t �[6���A�k+;b��pW?����Os8cIl�vl�c���T��W�5���e�M\Z���!�45a���^}İO��1�0 �J�/T�v��r��!�����N��<��Ԋ���	�|�{��q ���7��]���R?u@j	V����M"_*my���w�����Lo�H�o�P�����~�+�:���v�5�L�����m�O���ů�^hꉹ���*�h;�fz���.J^����;�Кt����%�����MPP�>�1\c�W۸P�=U���[xR�O[A��s�6^��w$�F�}cBx��}����,��P�t]��?0T
��Ͻ�� �[���g����8)|�o%)gc�C�_�11j���#�����u�P��=�����&u��y_ �MB���[��@2�1j���,+y�]����
�:,����g
���R�z��G��2��u�LiV��]�P�r7�6�S��R�hm o��3�'�'ȕ[D��)�" k���R��.T���B��V���V*��U��c�^����|�y~����Xñ�6YC�RzM+�3�Mj>x�w��B==~�F=�/6tyv�N�=%�O�zN�D���*4����P:�
z&zZ墮Q;���-�����d�F���s��[�u�LM��<;n��y,��_��MGJ����0_/;t^~ �D5��g�m��	/S*���2]�U��n����CL�5;f��u�³�=(4���B�Q�O���h#�lKv���o�q�#zhC���_���Jnc��������`�Qa������J �KZv���Ԣ��o��,�*�oc�Pz��@��J�|DEW���h�Ԏ�wM�fqbm	���)��hًc�Ml��Ǫ�X����*������G�i�T�ԩ�>�n�O��_�z�8T�Ӝ�.jjF�՜�C��؝��v�16-<$"��R��y�;��g��_m�2�d|�E�2?S��1}FGy����D3�F%���ˬ4�Z�~�Z�+���/�W �*7>�Ӹ��6����kNbfqs�æ�-�[) ���9�,
�(}o����c'����wc���9{$�=i[챷,��#jk�w��������A��JT˯� ��U�|����]�)�ؑ��g��w�ѭ�ڜԬ���V��fKJ��)A2%�*k�X��x�_�Ő��$,���W�1�t~Y3�2{Y�{Z����`��ZU�e��P�"m��:ʊ�B9r������P�r�X���LALa����C� !����z��~�V�ΡM�W�0���A�jx*7���ۢ�|b)~kkZ���R��u��,�#m�c�4]�q����#g��Oo�q@+gQ:d!K����]@���E�����܀M�n�[ �_T���9���ե�����ͧ(�Q��;�ޥx���{�5:���+C�E�/}ݲfbO��"�b�J�lF���D�OE�e�3��6��^U�vxD��4�te��0
%����,<�Y��0�UKq3�Zt/V��4C`��;�j�0'匩�.�`+i�Ph�t���P]�<����u��v�OX �fK����ȇ<~z׬Z�@}[�D�J�㪱�������&�&�����z���z73NZk̸���}��&/���2#oT(#�}Bb�#(���+�d\MNr1�٭ⳗ�7��?�9|/�\K.u��K [koj��n7�^���d�i>��4CG=����a��d����_MC�d�C�>��q=�?T��^=Xi�1�Ƃ�6�4e�M�p���u�I�X�ɗ���Ir�.���z��~T��\O,���rItR�l��5�mQ�|���>"���9�,N^�7��g�Lb�*� ͐p���ᴤ�G+�&�_��e���u���u�����h�X�mj�Z�<,[���d�wʂ���*i	�@�R5U,H�P�G�Gb��(�u�(�V�h�޸0J�q5��i\��:�R+�P���0v�/���w_�B���W0b
�c�� ������JZ������"e<ڤ�������2$":QNű��Y�y3w�W|>�ב�=s�r�b�j@���I�Q�������5-�P�Y�;`r�xw�d0���ٵ�@��'�x��*!�q?�w�CF�����z�k�B�[�`6v?3�Mq�DKW M�͉�c��7����"l��v������Xק��L��o2�F��*��Э��oq���{
���
��D��u�%ȓ�N�~־jp�Xm����px��'�&���mf�����br�v1������'�b��=�za�v�ci3�9�T��.�n˙��A��f
r�9zY�1��v6��S�ɔb�eB\�Pf����bi�GhF�f�E>wK�Y��lC��/�R)�@���-���"/:g6q����oG�o�m�"�L o4��"$���,y�uN�1L�j-�FN���gF��q�j�<�d�����tm��9�L����8:��L����?ܘ8�ů.���j��3y�j-��@��h�c�?<�%o�i�dxε��oi�� [���J����J-q�.2�"���~Kf�Y�ڒ���g<��ݐ�AC���ԃ�(�J?g�FչB&��j=.	�Qv{&������w�y)E`���@�!�4}���@.��q���wޱ�E�����@y���mP������K.�%=d��H��K?��M{�9z�c=�]�p1��r5� I�	�
���ʣ�OrA<�O/���iQJM�Q���W[-�Ņ\����.ַ a�e@KN���V�U�X�tP���pҬDU6�]���2�|�v��>�,{d<�͔�Ӎ�ݜ�zU8Ǆ�,vn��;F0~>�oOO�)/29�+>/ќ�׏�$X��ï#7x8]C��vb�1#�2W��U�J{ث{�} �=���k#RlוЎ���#��+�Y��+�����2݅��r=�M	��[Y>J3�y��VF����Q�:gGF;C,�R�l��1gy�J��N�B�)�"��<��h�
Lj�
����>�M\�ِ+�%Îז�'?f�Fl*Գ�,����.�c.r��*P����Q�o-����]D>���<i�����q^��}��$/��_�(?)���s?���Э�`�h�R̷w���WS�O��0m�Q�Q5p��DWR�J�����=QD�l/��y��ݍf�#�7"�9dc6���x����+��0��kس�t�wh}������i�x��k|K�	�r��'u��?��`����Y�R�ѐ���ƍ��'z��AI���o�|��~�M���N� /
��7�o��`Le��{���J�l���B�2e����˘tI��鲇�i2��o���~����$�6��4Ki2����)�k�k�DH �����_�^Z5ߋ�"@�+G"UNY�pS��L��l�-�O��j��I�_�C�W5����3���nֻ���41��O{�D�Y���mx�utsD[`�+`[����Ў5������@�,\@?��r;���Zdx�7�^[s?�M"XS����4��������w�g{��>�ќ��V o�2�\nq�YX���r5��5S��{�lڇ�໨�T%�C��S5wj��"�%o.�<��Z����iY@J�R�e����oQZ��L�E|�3$����d�bNа=��D��`؝*�:�w^��C�Z��N��AG�,f�y��(�,"��%.��v�|M|H]k��Ցz�EH�!��	QJ���bg�R�q���}2���(\��
V�o`�Rv���{�nX��ZX:�7�J�TL�Ds���������Jy) 'a���\��rQ��������4O�7If�:hrJ��~i(�t�W�����k&��)�s	�����%&heqtV�'������bb-ɍ�=��N��7���}w����k:=��A�a}YU�l��BtN����F3����lC�wDQy�8�� ���@����ewkr��,X�,;���.0������a����H�N�[��P
@�_=�$��=_���S���t�w{����Ng��;��գ�#}���9�@�<��j�>\,�ϐ͜�l�M���uL	o�P���9��E�p�6ƒ�U�P�kw�Av������A��ek�X���B����i���B����~�Җ�'�LK��7{����dc�O��~[4�c�`0�����e�i�_�>3�֥d��6|����g�Zi~�,�<�4\d'�Z*`غ���%�����y�#�}�+>}.�=8���~�Ѐ�#�?j�w��۶�+�L�c��dyp1W���U8�����<������A�i������A��@����V�B&�͎�����c�=Zh~���~��tB�w����zq^х���e�D�]�^ù!}{\R]�D}��93C��
mtO����P(D�/��ܤl��S��� +��W���ue<H&lڟmKČ#��C�J��(��,?i:��dj��s�5x�
��:���|�R	��0`�ֈ��|�rF�j��%6����Bn6{�dq$<؂���K���^Y����O��6{�\'M0jS��!P���Tr@�{q:��jԱ��R�����S�˄�[O2�,����X��r�F�^��>�A���.�[x$��:���&���e��=>RW��^_T8��૽��BB��^J1^
�n�C��y�ّ������l�eX5����|���M.����>�g
��I�dP�u��3����U�Z�:��i��6����߅��#N�K3�.�g���$�W�	�&���G��zU�c�dD)��>��Ad�wH���D����zc�M�¨��T�Z�<p ��(���{Ǧ1����!ۢ'_h�.(gd�:J}׀e���4d��:�'���)�f�B��qd��XR��Q]@��r%���F,��w�=��.l�uDKً�IG?P�^xjY6���c�3j,�ɗ=!���9����k6��R �CDR������֚�^���d��a��~�M�;%$�\u/QIm��6�#��u�����4�Y�mq~��PQu�`�I [@�v�g�QC\p�F~��-�3<���%��u���]�4>,:�&>� *>�˄�_IA�2�����`խݘF 
ͤ�mb'a�3N��\����(���QAn�˖��@�V�dD����D�@ΐQ�v%�E���phm�O��#�Ȝxk<s״Ɛw��ǚex|��yI"5>1C�j�2͗�E)��]��l���(SK���Q��V:�ˠ�<��cQL9h ��'�m��R�G��P���x�}�N:#>�3{T9��(�Ij��Y�p��߭���BR|<�p���_L�y>~�R���@7lZ�jE�K^�Y���Ѯ&���Z�Ӻ�9
���{i��`M0��_�z���v5]tl��E
?8���xR� �d?[�,1��������.�5�����9��䟬��y�vU�Ȑ�����t������_\�6lR�^??�~������1�L���>�S��]9�X��В5������+V�cA3.~>$���7X�c	eV������įI�J��!��EB١G�Ԡ��f-X%����3�|~������<*E�ڦqv����������^]�L�\����P����N�U�v��m�
���cZבҜ*��pw����4m��y�r�ϒ^���*����Aot�(q*�72Q*��pI�/�"�՘���V�\��,X�,a�\�+���8��4�f:B�2Y��D�w̭]�u���OAWܰ����l ؠ�¤�!���Pt��#r*=��2�&���(��ߓ�U}@��?��X�'Z$g�9�T}�DP�P��>Nނ�N��=�4�׉��C�2X�$�vc+���J�z1���p�+�s��3���x�D�3���"8b�5rI�4�h�.Q�d:h�>#�}[���(����n�����(���{��;���0yh�m�q4Tcw�X;cT4���2�5�M;���E��p�v�����'���;��ԟ@R/�
n��8��e� π0��d�jGY�z�������(�՛#�Pk���sQ���^�չ$��ܦhd��n���= �h!_̺�ovxYȮ�g��ꉛ7�;��(�͈^���W�m���*�V��{&��9;��-,>�qN#����Ź9I��()����xOiQ�E����Bo�w��v�ۏ14�]��,;ˉ���E'\<���b�ns���C����q�*���9�z�S�B��#��1�E�zá��+il[����}�'�&�s��/�w�}A8�`�J�:C�S���)u��A#I�1P=&�z��ت@�'����YP��}=�[/��s��S��f���In(��5C�������3�m
�����s=�.�Nіѕ���o��+? �q���`� ]�����Q޼�8�4G�ê� ��z�X��$1��1��5ffgv�����V�B��b���tFv�h�㍋] j��k;����;O7�&��UI�*���Kɵ2G1S�ԭ}JBNB����d~�����XN!ơ7o��w��\�p����O~�2�Ų�H�W�cd�A�+O$����Ge0h;d��ۗR$�d%o� /�6�5c�K�$~,��Kn\v�T߇?�R:\�ڵ40@|�,̇�I�ܻ�$���e���r�:��C�������1��-��~^]T�W�#=��N�.�I��ю�?&3^A��;n����1O��k5�����'�$�h�������~��5g$6��ʁW�Cm�k�J ~$Z�o��~?�y}
`���o���j!��:�h�&Ȏ�A�va�Ͳ������w���y��U�A�����2
��O�6K���G�7/�n{�F�^�X���Q�^��ƾ����8^����o���ê�3���~��x�V�&vg��;kG�	��cw�H���ڡ�T��nf�ص����I���B���3#?�B��U1iq�&wQ�=CU(�����3��
"Ӓ��@N;1���D��d�ɢcG�� �Mi,��_�] �U�V���IΞ����HIU�_ ��ŠNk̤��H���Qȉ��}�E���̘�)?�� �>7D�E{��lJȊTI�Α��8�t,�X�d� �0���ګT���v���������g+1��M/�E=
�N�SLW>��P�ɇ�>zR��2�`��_�
��;��8.���C����p�t���1"��"���e��J���*d��R=y�}h�y�R��  �ht����4�j{w�V��~����қb��?�-�|+9�^p6 ��D�g�͘���'s��;�N_�nk��,��4w�A��3�GwW6�K����bz鱺Ur����J�UFN���io-�Į�/'h�A:`�ҩtfx��o�U�5�������������1w���:����Hf(p
((�եr ��F�kv�����i,e��_k9�{�j7�g�����qEA��_�$+d�����#����f`�WlN��dp�yk�\�t�s���[��W�5�ZG���V}h�)�z	�_�Z{�r�@���d�����䭮�˞�h|�q��D�v�3��0�vZ�6��p����/3�>U��0�L��E'?�2Qd!�ӁH��A��c�R��/S�/�=�@����H~7�/�&�~�cKC�S)s	ȷbI{�>�-�Z��{;Ж�X|t	`A��uZ&�PU���9d��Θ�&�=�T�s<�����qd�e��uN�(��k�Q_M�Q}W�pU���F�Y����i�o��ӂ7��@��;���$g�����,�&��w~����B�(L*��U� y��ʉ��E;p��Eu)�=����U�u��ڗ�^\W%:6QQ2���a����z0����,��`�k�ᝑ�b��<���&PȤ *!��)u�)�'�(�����^���I�{�����	-�94�:<T��W�>P��I���M���u,�Bz�MtHע4�F�͒B�U$���%m�q�w�Tb_���t����/%���$�D@{�P��c(1p�����R)�/�F��2=xz����\B�n��C�i����l�k��R�)�Y�Ø�K-��`�G-�.�2/�����v�旄7��5�Q��3�D�S��~8���&P����2<x�Q�!��4�=�>g���=xʈD�j�@X%�u͙W�}�����Ta�μ#c&&��(�o��V��\�U������Z�\�^�#��4ᒧP 3�31�p�ᩩ�OO#S��:�ə�,|B	F���}*6��KV��Zf�!��"�q���k�~�*�`��,V�P��pv>��E���24��
�\}�G����iֻ�eD� [��a��ڻ��E
)�P\ӁK�b�YE�D @�)�oS���v�b�$_/�y0��7BrW���҆�8�U��8��#x1lS���!Ǧ�O
�@!M0M>Tz[Lz�b]X�$ξӓ)�9��o��j��;�	��.s*~0=3��3�Q�{�o��%9���H�UVX��_�0ؽ��߷�!5]'s����ӼA��,�i�iY�^&��J�#��G��>����F�V�ݰ'�胀�fG��[sF݀Ww6��P����R�q�5dD�����P��3��ϓ��c�;�V��q��}�B��`�W�{��1����xtG�HA㥧�߽���v{�\"�19�&���0��u���K��3�+��mF��k�RPW�o*�=�v��6�s�9��f��?�V�����y�;%��]Fn}\��\Y�������tD�t.��c�HY�XYds�r�2�_#�U*��o9�G@�V/��r=��	CzU�A7d=T�ًXߒ�Y
�:l���-,<�D��TR;�Et���	��ձ1���{Zi"+�&4��ڢ�(�2b�[D�����/��G^�%�8�ڣ���r]=Y��(�)ʃ&�o�f3��̼L�����0)>�4�?7�/׳��a��ŗ[`�/�Z%��bQ))D5<�GL�o�gNڮڇ�;lUvz/ɷl�$cp#ㅟK�p�=�[����Q=Zӹ�G���u�-!ۻ���zh�e�Cu��"/���=̛7�I����kL���)��`���#�b��P>�$P�1!%���Xp�C�Y$��z���˴����-m=4��t��ٓ�nY>����f��:f�Q�r���6H_�Qk"�����^(C�p-X�D��<��p���}���K�i����/*#���r�{Y	7�$�y�2�|�e1�3��+��d���{ ��|oN�5��B)*��dii� ��	h�ש�G)��­��ʰ�Bu>� @K�4@��J:k.�yԙHϩɑF�oP�z��� ��Dx�ڔX e5���\�͝8�|J�V�� )�A���l�|K �D�وQWo���k������1U�*�}�ҕ❖�ߓ�� T,:r����$dq�c��1��>PӵlZ�=�m"7M�*�)i+R(R�d�â���0��M��E��y2��p��V�x�֛��A��L~#��"W�cށ
�l߅_�_].���|���j�}1s����=v;����};8�^.��?��z�"y �\�CW���6�/���jB@����k0j=�D	U�tW�#��f����;��^��!ԓn�h�/��,��x��S�^Dx�{�5������>Z�����������%o�@e�j�\�95>��NJ��J`���.{K��
Po�ũ��,b
���*���Q��H�4<�$�����ת�G��N#�:���'�/����U��&�������h���ϒOP�D���w���n*�vo������� j����	-���I]�����	����ɲ>��J��.pB�%C����72�����ف��JJ�b����5�
�B�^��ĭc�~u������[�͔�t-W6-��"�]�n�`)��m��ű��\��@��䲋 �?��}�z��zn\�-0�s�c5��$�c�k��0���t�*�ޒ��|=a�ȫ��;0	��UZ��P�$!y[ku�\���ۈ�����١�ay�Z�@$����E��ͬ�ف���Y�f�� ����ZD�~�QD-�d����D��K=�n+����i��9�>*s�b�h�
`'��d�> ��Q���gm�/��5"��;�U��qㇵ��A��<2H��b�g�"�M})�*J��$HhK�8
1��b]Z+���g�9�&�G9 ���0!_Ny�!j:>A�/F�E)�S�)�-l>t�S�����[g(U7�*˒�P�˄h`�:�)��T
�Q�fn��W(�k�&y�6�^O�����H�S��.�A�W-�>r&2mx��i�S��d5Q�X`�ɷPRѕKG4�=MȠ�*������M�Q�~�'��h���Q%�mE����<<��`���e}G!�VEkFA�d�9f��� �3��@��ܨl�� J@��*��6S����;���i��џ�L�+<oi�F��~�ofUٺ�8��W���-�c�h�X�9��ym	�<�nlᏥ�N�n~u4����$dژ��,����W�;
��.��,I��[�mu.��s���?t���K�	b)�u�^�9~|�ė��r�ʃ:�����CS��'X�f��^{�'��4O�`�Y�l�H�4yΊF��^��(+q�j^�A�(5.
��U��.\&<E�c�ˢ �G�\�p���Ro�N.=� �B(��m�h#l��O�T�1�nKx�M��d�싪Z�x��lv�%_
�.��\5dqJ6e��'�#�3�S,�j�!�7��P@N�5�
��~˾k�D�X䧚���h�VC�gE��W�+I�����Evq��Bga�7�r򡳞���5��tm��1�!d^S�{�]Ы�a�<C�;��#�_���q(Y�<tA�'vpo���U�1#�-KJ�5��FS�q��st��$���ˉ�����x�-����Q�h��DѪ��aڪ)�uT��0*6��5JE�9�����,�Q����%�-%T���!b�D��8<��S�ޝ-y+�X�cC���x�X��7�Ȑ<˕MpP�嶗��II�s�8z��A���0ǐ�,G���m�X_e-����2n?�����S�FR�l˫��U�)!�r`�#���؁"4;p:ӱ��0 yn�n�,C5|Y�{�m~G�p���J���V}��`�;Ժ���9�������hL|O�T̤T܉�����#E�v�P~c7_��r�Q�ꁏ�%�����E��|��e�w�~�e珁-�-[V�8�;�޶�!����(;�����+H�^�v��?���Y�����AUJq�h�rGJʹ��M-9@a�衤���Ͷ��y3 �����RH`u�����̽~��N���:�G��c����y��H{��'O�[>J�ؼ,[�en0��G���w��s����;Jc�Ꞓ�˪�Ғ�4<�T�z��H��qמ����oV����CJq��_���$�X���T�t	����k�[��Z�4�0=�H}��ju��U�94���-����������(� ��v��P�,�g̊_w���+\O�7����ã��wLZb���8d0ԘM�`$˝��Tk[y#�4�� �������R�O�]+�U�8�\��<�:H>+]L��Cb�����S�U�LXaɝ��/t��p�&Q�W��!is�`�8�
�IX.r�����1]~��D��,|�#��`���&���Sp�>��Ar�����u������-k���ֿ�߽LK���f�S�p�����'qCv�Z����^��4�&Cvcf�߽�-_>R�+���ʎVE�ѽ�}�([�f���N��B��H��g�R��=�EʚI�
F0�@�7�G��]i<%ܺ�s�z�ڤ5eޣpx��(n/�U@����=�j��ܦ�C���զ���U�:E:Ц8rF���h�v�";o�6X�Z����������dY�͗^��-M�bпĴ s:�1%z�����Rpv�N��x�wF�����mL�o?@��E|#�؛!�C�y�H(��<��Ń�@c�;�����7U�<@2ށ];&�O���p2�<�mE�,+N�C� ���:��Ԡ>s8�V�['�a�H�#/�
hB�h&h۱j^�����7���8i��������:[:��BԵH��Ք������()L4���ؤ\N��`�{����e����>�����p6��HA�LE��#g�j�������t��
����W��;��(��o~Yٽ[q�<V~�i-�q���0�{|�ϙpb��w`n��{�yw���Qe�o��#z�>T�xz+��׮�������W�Y3u�Lk�cߴ.Ҹ�Z�"dA�|�#�1m/J�I��g+_�i�KJ����<h�.Fӹ����3�5FM�r>�O��ͯ�����JJl&���3ٖچ��梵�^r�}l���Y��#�.`����^�	�T�s���d���g�w\{�Ku�pbN�d2|OhۤM7�]��W�������m}FL�(�e��a���s���w?��.b�tKն�OA�����ogO�О�����1��b�c[xK?5�^\Z5���BL@11��Ѓ֕��,���xiƓP��D�b��	/�DYv���x��RO��v'����{��=�h�!����-�xp��k�F�;Ϻ^�}�".�t'ı���hQk�CQz��j�xi4��H��߰-=���#u^�.٘x��΂�H� p!5��Z�P��:�RTW�TYi��KN'O�ƛe��*�Ӹ��gy�q����j]uqox�P[� ���hf�pp l(f�ut�˿5U`�40�"_ӣ�f���K��1��O#N��x�ˠ t^��wL�F��%�[�p���+щ�]F߶<!���Q(^��-{-k���U��#��a�A暽`qR��t�c_5z����'!R��BI��6��{D�S����`���ky)C���|��N�;�-@A�-T��_෌��y�J�L�&C� �X������[O�G,%$�0�M+�	1�Ǥ��̬E�ߎſ�������ᓠ�/K	M��[Ӑ=B�l�
�JEC�
�0X�p�w}4b��kftR�0��)��K�=�?l�ڤ��p��S��SZ�HEX��"�J˼�-h�^��+dk��#z~�#��I��mH��y~���ـKi�}z��pɉ3v��HT�(�~]�!�R ���jz#�B=E~~��L=�?�������*��|�ոrV0�ֿ��TA%��6_b|�M1���]�P�;���[��Zò��ҥ��r��j��	;�~�c�jl�A�a�U�(y�yc��=���`:�t�ߊ� �B��(ASO�,j¢CC���fD�{�B�w��cK�S�����}��E�s<�{�rݯ1cR�7�vA@�T,)ÄYbC���V��v(��awI�C�UaCTc"xUN|��*�|�� ���y�� ��
SЀ���e���0���x�����  �g%℘�<���3���P�M�t{�Ν�� �,;��(b������-*��-�-ũ{��SY�Z��[�״^d���|�{(�"�+�(�@B�N'Uj��v��um{PghK�iwq��&�����p��,!�8q��^^ܦT���Q�� 3S��r���>��H`�A%��~o�Cc�5��;�V��h�~m��jz5���B�r�9����2�z��m��W/}e8�j��������:AVF��8��=���AǍ�auX�R�V�0�\����?��J L>���1M9�l�Q����s�	N��N�8pp�,��[@g+C��ف�9���"�CG6��*d1&An��I&f�2�ɅN7�xH׃��j�q6(46d%��S�r�� � J.?��G�9^� �Y|�.���6�?��n�˲ƥGj�"�����Bh~V����0D���U� �y3��h���s��(S8��f=}n���R�}��E�(�t^�C��H��;k��p��ܽ(X���՘FR���ꗾY�����YNיtD�nn�� ���~��T����z�'�U��$E��B wg% �G��c~t�T�6	Ԙ} A�z�B�F�j^*��$�)v���O��-R2���I�?=��x���������#�ˡ��4��{�����+��A}tS�.ϚU�K~��q�(�A�W��m]� �ژ{Ǭ��^Ɯ�)˃���wf��O
v{?�������""����e�F�H�hY��D/ֻm3��!0�6��&�� ��>:�6�0.��k~���^�
���n�H��Zz��(�ˌ���G�{W�Oe���R���vP��7�)@�l�W��҉���2_%N�>�}S��V�}��2��(�dteSY�_�ՙ���X�4��tG�!6����<���چJ-��A�j�H��i��� .�wY�#;2��'Dz&��
�EO:j���RiA���a�~Z�\sR�ץOt��-�/���1��rU���<��o�"/��'�mr��m}�L�h.u�����D��J�By�l�&V��m��I�w���(<��C��	�e!�>�c]�@4���3��>|��lja*��ʦ�x��KPd��X�y�4��73�=od4��c0��?~cG{B�Y�T�9ҡ�g��Hک�V���mƿ��8A}I�� ����Ph�B��#i.N�!�����b�3Prh��m�t�e����::���H��ͬ��,ނ�\��(�:Y��|ۍ4h��rȃMgp��4�-��;E��TE[�osjO�Q�l_�uhά�ƖӴ��M�Q������k�uav?� �	.]cP���a7�mz��ؐ�ZX��2���>j��E��^u�?��@m_ǻ��G�I��_�aӭ�gi�=,Zx�!�"h�� ��"��4tI:��z����b�-�'�4�|[I�����a�(�%&0�0ߎ��$貙?�g�����Z��y/�|@_�v��vvE�������<\4J |�3_z)TK#;�����ڥX>l�>B��k>�\X��l���M�����5&�/5~pe��>@``-�g7j�#��iFi�Dd���9�, ��M��<T�ΐ�>�/�P5�T�u�m�Ԓu�9l���%��޴Q�\P-����2��9FT��2H�ō>	�U�W ��A�h�*Kv/%4\�RI�@��9�!�B����k�C����/��B���{���
���7�IiV��9m���,������=c]A��z�ha��?�%�X��%A��=��^����w���H�N^�!�n�� F�}�5Fw<e�*���X�x����H�y������bI��=M�vP�`���v<Js�{s�ml��K�d�A�H#�u�bT����-�hJ���e���;�$�����y��8�C��g��aC?��<�J/��걹&i���m�d���p����z�w�o���	 �IK�+��ѿ9U����֛턍����c+n�>p����]<?��c��b'�Z�󦔦�-t.?/�5A��0���J��MW�~.1�N 6
|�
�C�1"�7q���9��\^q,W��?n��ى+�"1/�?�0/��䎟�3�j(I�=��y�t\���"Dv��BjM���}xk��"[�	��m(ha��ўV��:�C0����k-Ĝ%'m)Kwxt|���������˿Tr�P�p�Hm7���K��y]����A�i��j����K���RB�	�B�$�މ�|����$����g
__����bk*~�g�\l��6:�d��!T#�Hz;1k���ok,� �33S-?R�3]�	t�XU`я���?V����#��U-���04��kx�J�Pr7߫�[,%Sa�#Q&Si�A<N����X�N�T�R��i�lA�jx���^	�K��%�@�i�����k�t2��@��Q�&�f��f�]1�'?��N���R����y�e(N�w�l�������1����=.�έ�����\��7�������l����/N���[f5��$|gL��5Z�1�����^�6�M��� O��#�>�S:����T�޵@v���7Z�.?�J�Vd\F����\�~/ԉ-=a�Aq�Ο�V/�HhWM��	��Z��[d�R��y�u��sQ�!��BK��
�H�fޔFsQ�6��{�d�� 3j�Oi1��m��f�)��q�X�wt6@�E�@"�IDI�r��|�\�u�)���r�o��>s.���&B�0��И���f���l)A��K���0���V��rmBFF��&��Z���<(~�CE��#���������7�8����T~��E��R|C�;��q�5���#�WvdOW�D��GO3�O�ܱ�38x��7)t2l�>��':X%��X@=<�4��^?������ܟz�R��G��s�;zkA�.'G.
�V��1����N!��]���޶�z��
��Z{��-N��]TuhH
Y���m�ѐ�w!D2I6�^4����:��i�|�u�s����C3A[N��϶h5MA2��ߚ�*����v�oEj��-�	�%��TWfw}�0}�ԭ�!�%=��5�K y�bSq5�zlY��_��W�V��|3p��7Fz�21)���E{��%FMQ�;ؠ��C�2����<�ׯ�,�-�<�����f*�2[Ӫ�����ѽ��� �� k�8�ݧ�aq���^lR!�v�zz�b+z�EV����"Wp�����\D�F����unR�A_<(V:�M�(�Xў_�Ԥ���ࠛS���9N�n���I��L��N�o''�q\a�
m�H(�������F��%�Z����ﯷ��[�y =A��[;9j�6��7��5c��������4�2�Wk��ͅe��}5�P�����Q�cY�.���u�SR7�&r�v��8�Fk�ȗ�/_�y���5=�F�
��@�˒���
s��O��;e[�������ӆ��W|�Y�u2�j3P|E���x�7�|���!�I?�����:�2�Y�n^+�0�+πQ�(i��ԱǇ��c���9m�T/�Aia�Y	[�ϊ�oe���N�����r@v`n~��A�#��$�xC�|hƆe���ۆ��?lg-�X�b�y(����B��TWߎ��~F����Qs���aVb��AayBy�G{��L�~d�a|QH\OPmlpx�>r�������F�=��V���^�|M�o��C���m ��D��]^�瑚@~�Z��j,�WM��[��9QRIܧMPG�9���[_$�ݚ���*�����x,�ݺ�:�Iw��c��� �	���iج��˪�]���\m��)t��|6$"nt�5�̀ם۽�%8�<Fݑ�
H�[�r\fs�E��<�`�V+C��d�j"G�5�+�\f6txυ!��S~�nos��9l����xa�F�����&��S�Y�Ϸ^Ym~�ރ���20��a�3?�G9��9	`�Ԥ��A8��yU���XTG�{�M���+�s�/&���WM���r����jP�>�SE�鞟�Z����V��D���Kܝ�*h�f6q4#��zK ��|���%�h�irXH/a���dSu���2
�(�p
������ ^��M�-��Ҏ�5����
&�`8�U��?��:H��d��Y����?���y�Z)Ԃp����� vSW��;!
�c#��q�����A����ex7�ٻ�Ǖ5����A#(>���XM��h�b�t5Y�eb�i�R3О�yV�Ӑ\��1C�ht~�������\�Yu��c�s;��Z��6�� ����%�}��eK�v���F�<�
�=Vb���>*��ԣ9��ǧ���`����n'�Q�� ��e�^����%sצrWF�	�%?��p�E�Ae�w-Em�d�-w��J�*���&�Wm�(�=;�t20	��<$=���I�t�1}�Qj�,�Ǖ��+���"�?B��J6G�G�*^�w�K6��46��%�y��]<s%�����0\�*QB*�N�,���!h���:�4�N���=g��Hf�,����K��o� <|�L�(6g�7NQ�>\#��J�	��$��s�sn"�(�K����b�K��T��t�d�(/���<9���v���Y&
A?��
�����銚�tl�uW6F�A-��w���`m�_��?lٸ���0�(m��!��q���Y�����M�tG��q�����rb삎mj�kp3K1��K;�'�5���ybJ���4�R�] �g��i�-�<�v����	I��r��؃��Ұ�F��e��a���*%r��.��X)��f�|�bM?h��|0�voH~U*��j���si�����z��#l�}�O��"��9X��s} ��1�^���%B�!�3K��*}D+��l8)�;K&�,�P��L�>�۹����S���~=0���9�Q&5\�]� ����0�G]��!\W7_��Q���b�	��ZN�7��`%�cO�#zڼi��0�`�N\מ�rk)ֆ�ʀMP*)����8��т4�|Ɉ9^�&Nw���a3���#�(��M٤P
t�<
Ic�h��ɮ%;�@�$<��ArtO�,��cl3�&�7hk#|��ضq��}��qjl/�zG0ne(��5����D����5�,8��z�	z�"��-7,�0Tt�[�M��`�����ϴ�~v�K:]w�>3F%Wo<q���i�	.��t�9�)�e��.@`Z%N�_Xu5N;w�s#Ӫ�?!Q��;�!bbN�=vW��*�̊�q��ݦm��"�s~��p�a\�� �x�\�arNL��{�a����Zx��h�K��"hI����f�<��`������������>|�@���I �.���u���$�o��i���i�I?�"���>��K%�to���D����\����Cu�$�!
(�T�p�`n}j��p?���ԁ�I�<s�,�{<I|���P�ޫYzt�3����B��@U'�`�؂�ny�͜�� ������}rl��콥��e�y�ף�<`G��ls��j�vyć��E���6G�S�&􀥧�/[l;�����	�ם���qq�H�jR�%�9���@��
�(��7Ё�p���a08�S4^�|�K^i��K0�Z+ �����R�-��ƾ �=�K��� ܏�����ߧF#Ӗ���p�⋛^�b�0M�<�3<�L�"�FG��)�i}�����8W�9kH�2N� 3��P#˂NW(�Qɱ:�@y=UIh�6W�y�9_��臲#���.������w7d��߷X*���������}P�p'�]��&@k��A\���U�j�q^��w�3�V(�3`�L��c��p�F� O����8�1�l���z)���v��;+-�0�N9'#{�ק�\�e����4��Z��\�K��~���h{ڷGXd�z�cuG�F����� ��* �a�$?v���vD��ː��5����_O=.�V�-�����f��c�VA�f��x�qc�֨���0�N�J��ޅ�}S1�?��!��g�I	}h����7Nm�b,)�Lr�ӓ�"DZ��YN=h�6�{4��g��	�)[Y�,d�(
=NU�C�<W�0I�g=���'�*��Ng�}�*oX�e�o�ޓ�Z� �6�T��K�,%�4�Uf'��]x���	8	Q�`��}�^�1{鏪	G7��Y�x� ��#3XQk�'a���5�!S��*D%uV�2M�VȞ4�E�4���H#���@-fb`��R�t�T�и ��-e꠾��U� x��K
�&y+4e+g˗�L�:� o�χO���۵vp�h�܂,[&��5�Te��e������e?4.w�ʐ����%���:�hCGW�����I(��� �8J���8X�ǀumE��z@�k�x|��#`���.��:��]�&_��Q��y�-E�+>Qk���j�W�f5d) )���,i�,h�;��a�h�b�W���%�n�jb��#��I��M�c(�o(/�gAm͐�T;;�a���c��Y�li{�ӝ���ô�:�K3�j��x�v�DВ�h�w|�e?�2JҞ &(��`X���)���2�2�v���n����t!���͑S���緐-pϓk�~90��dDH�����L ����L�Vo�2u+"l�f.g�����WAG.�hYkT ��>�&/�?rM��$J,3@���o��Xp}0�;��`�X�R�]x|h�d V�93�A��#Zƌ�Y��R֚�!'�fR�|J�V�:Nf�OPDiU�p0|��m_��_[R�����Yъ%�(�al��N��;*�=���,�e��b�J��T��ib1�ݲ/Y�k�_�g��]��
���6������8רxk�bm5`it�k���E���m�YȔ�>��'�\%�{��UP=���_9�O���r2���"�����Y��7�?��$-�'�^`�]QD�8.�5"��nu�OVyȚ	���;?B9QE�?w�{z�(�\��9��.L�+��4g�,�P�;�5O��$X7U{]�<'�_%i,�1�����mߑ�5L��B� w�(��?)ͩv����4+U~<N�����UA�Yz�4Y����t������+�}V#í�K�њfU%�!��"nW\n�	�e]w�/�޾w��k���Пagn^N�m̢�ŏ�e��t��AQ���%�e���#?��e�܋�zA)v�Ʈ���wEЊ����Lf$��?����������JS�����#"b$.}�I7e9褍ǲ<������&����P_K7�,
�����2	[x&k�'r��n���X``��Z�
��F�ߧt��Se�y��NZm�@���ݨ*84֓�$��*�%���9�]�S�" ��3	Y��L��e3ń�o���p�e����f'���wz��6��N"�񭏁�������2��2�����_���^��/�w&O���.7��8��E��:��ޠ��O<�Th-�S	��æ�+�w[�k��,��8��$��d<��#b�i��d��/�o�<_{�$�X�^:"� �T����=NvN�*��lƁZ������o>H�5ݮ�̕؎I�VEu3N'Q�׋Hu�ݢ�����!lpSҁ�K	i�����N���I��G�(+@
�#n�q��2��Cj{j-(��A�d� �c�!�#Z������r�qg�28F�[˽z�و@�ӗ�(�?)�r�1�궽E�d2\������ö��P>f��� )G���>3���m	)�.��#g8�0xH8���0��陮y���8��!K/M��ٲ��	���tVV �O�H�͘�w+�h�7���/]֯g:,U��H|>x���,�C{f�x�]����B�fU�H�{���R�5^<Ph���P%FfC��C��`��޵57hU�G�c<���ѾB�'벖z�pBݧѳN�Ø�<|:�˴�� cb�?U-�=�1��,>,���iZ^|$c��
���hG�D��	��-�VćC���hF�"q�6�����1*N(��u�F�nMn>�#lȭ�R��6z�08�i�?:	�P$�p��ܣQ�sPl�W�[<e�[D�Ea�T_��N��K��������Z�J���^�Nb��Y?�K�3�Y���W#*��U���NhL�C�q_�6�&�c��,a�X�51�Pr2FvQ72�Ŵ��-�T%�/B��ej�.$��9j�5��6	@�ˋj�l�q�d���T>t�")^��Ir�Q3���6e0�6-�?K��-�%qv@%b)Z%�TW��UH'?���C_w��s�]�0-�5C~hm.Q���uQ���_��#��4���$C)m܉E�B�Z0ҷ~�_�x�;��oj/`��U�R��,q>�f�A��4
��W�E(#��A�q]�lOiw{1&ɦ��9����U攆Ĳ�]rE��S]!�{'F�(����y��$K3�_$q{�> i�-�a��U�����az����_�˲���cM#��K�ڌ��X�A���0:��=IN����!w5uoS����§�V," f�	�IZh�u�
<�5L�����A7�&?�B���ϸS�o��:{��z����?��c�E(��z��<$,͊�d5���}��[=<��W�q����ت���vI��mC�e�D�w���S�;��虆d�%� "f;����Un����)xZn��϶��{~w���.իxVa��F�;F�-�v���XP�q���?Q�9J�.!�ن]?��|��;���<��yeyJ1��k��>c�=�ש��
��ع����ؐ��Y���P:|}6g���u�I�N�h�ؖ�}�K'}~t��a���Xxx���<���mO���U.oп��v���;ˎ����X���gƗkzb��׎͘6��S��0��k��}�L��!�{i�&uO4!�ң=.1*>���@d]�s�w$���~Δ��B(��y[Q�aݚzp�=�)�{��3]֋�7M9��dp���n[��{o
���Ba/��X��|�֐>�EAR$V�MdfE�w����h"���¢���ޠnp{W8�/d�Ȉ���d��r��M��n(Z���cm��Q�b�	d�P��2|d�P&��(�!\P���,�Q�E�����nպY�$�0�W\K����:���.A�}�������0�ۯQ1��'�O���H��P���qL�º�$�n�+�uk�ZQ:zd͑��i-=�x���l߉�%k�s׈� }�xu���J+���/��~���X��:M������ȓ�)��"ز6����yMyXґ@�3�y�\�l�D� �*��	��Pގ��{�#3�~��	a$�������)���ړ��<U�
K[�na�a���)�q�W~>�	�/�"Λ�JڎoʪMY:�ʴu�Lg�J�]»,}�̨��n��º�!�ȑfFbaw9�u�z��\���<�+� 4j�#4�Կm�b,��|s�B�����ֻG�{�^�53�7ݛ�'�	J����Xơ�E��/W-��I<2�k0΍���D���:��S���C���E|��e����՚v#%�	K. ��3����iН��퀴v�M�9cXӻ�5���^���JRJ	��x\�l	*P��Ĩ�g��n��#vO�#̼��X�t�1-Iv�%J�b���<����%�`�聱�Q���J�(Ǚ�0҄��ߙ�)i�uQGR�?O"��_�Ie�cE�����ɝ2ĈN���*�o�sY-$���������E�Pt�����<+5����N�+��*��j��J��B=QA�ؘ�u̗U&w�����w�%O��D��Ap<8;\zAUA��	gE2V�;[��[�R�N".�" ��T/�����Dy������K�0�BQ���87~�j�L��_�`�X��6_M���@���3;�sJ�Λ��z|t>2��̀�I�O�f���V��[QtBdM���E���&����,���f�Vg�CΖ��>q56� �S=Ss�Y��w��*��\:<��z~>�N�Ԉ�3���u�R�-�����u2Гx�݉�kE|$ù	IM�$�E���
��O���lg�:�Hf��F��ւ�z/r��ү�p���m�m�������rTк"�f�|���)aZ��13��ih��=l��7w2�u�RD�����������Lr@�����ZGѶ�x�}gp1��Y�i!7D��"<��u�})A�;��ב��V�X�����`H�.1��	[J�'��@�mD.�<����߆��$�Y6\�0F�#Fa41[���!~�i��&�e�� �O�lr�9��2�~j��>�I����m:�a�o�Vq��G7��q��]���@3�9P��auO����?����˲av��S�wĂ���Ii��e��b]\�;�l �ь|`�'��K��7FvXũUpg.�P�	����d�`�0���Oq�VA�ݼ�GG�3j���q��\7����ko���>Z��OC�z}
X�Zͱ�o�ך����GZ�D\;�?�n�A����v�;)@RH#^�,��E�M4�TH?s+��u���z�\˙���x+5�Z.Bܘ�F�nc`6�Wlq�^��T�e��O��E��t�p��G�a���ֵ#B�Z�A�o�u����J_F���Mk0-`��_t�F;;�c/����M#�8��#�n��tS�*"xu�~��^ǎ�|U���JFk���*f��U��	�H�w�T���t�Q?ހn)�&�;4����J���<0���0�k�<TA�x �%r��D��mRp;e����4X+0��*S%*p�]��ۿ�\F���/�u-��a8Դ�ZI��BJ�s��#0�_�4�:��E'&Ƥ�n�Ay�6o��M�Pxb�C���/?��\,}b�*�0�Z� ��
�LPB��{�@Vd\���#�ǃ���m���n�z>Dw=_wg��;�6�C�1͍��1�`��4۩���'& X��V���w�s�7��܇���O�@G�P�7��DՑ]Qmdp��)������௬.<���jk�S7M�o��E����{��r��s�p�Ͽ����5���D�$��m��M��=��=�N�.XՉ��Ə� �`*���ɉ�:�.��$o	e�Y���b�̤�M��眬EFRZ��4��r�k��Oi�1pv~�D���+��Rg���=#o��0�Y�r
�;���E�� �F�6F�)���ԣӳl�� �=�v�*R�Ղ��f�T�M6���7B�:�ȟ�?�;g�ڜ������w:e�NP�-��\`�!���Pg��ULE=o��/�\����T�4\�+n�+�t�U"Γc�y����J�e}��D<�ǿ7=������Ě\�*f�F�#<����,��,�#��s��^I�����9 �v�Z>\f�����������b9���vZ��?�4�'ǎD��pL	��X-������!&s�׋)4W��?����7AxO���5�Sb���`�F��u�$$)� H�/_�O�VO��/�{���N��g�EN�����5�Ӧu).9��B��k=�T��߰�P]u��l�˂�}�ួ�0(�X�i��6����ɚ��n/䩶�_�L������q/$��Г�;�|7|�ĭlN����y����/{�������ɞ ��(�@���S�|����*�	�ͮ��k���.�8�*4�W/f}e��k�U�g�z��jٽԙ/<dk�z+]�;s(g�{�1���,����1ڍ�Ꮤ9�ʂ����_����q�䗽O�ʛ}�m�9\�h�E<y���-��mܫ�q� 1��&v5 �d�V�,�����V���o�={�T�����u���������38���D_H�֞`X��|-�	m>i�Y����p��6�5D�\�o)�xѶ\���xP]�@%:�|%�g���Rf���y�Yej���i�15�
,�T�n�!����{B>0*���Eif�i�%Y0ߘ�	P�X��W$�9`ݦ�ۏ��9�:*�\MR-�~���}ݧ�.���"���*��}@�p_4p�t����Q�W#��O	iW�E�� ����&��F7�(1ZXp:�bX0ٞ���l�,����e�1��d�x��mvt������D���`������>J N�@1Y�nF@"�5�����O���f��E� �qc>�-o��#`�Q���r>ÜE-��Ŵ�tw�'HQ�J"씔�Oa�΀�Xx�3vP�#�e�9FP�O+0F�N�{��K�f��1!���>�0~��e�IW<�ئ\I,l���Rs�̬hGLj��s
>	�m��A����KLZ��62�s�ȳ|ߓN�(���41���%C��]|�s�^�i�*���{��8^�������,�;w`G�fٹ`��=jO�НPur3ޗ�	�t�w�ͯ�c�?��d���&Z+Un`m� {$T��p��	w؊�`L����Z��o4IHޡ���a��m@?�M��x'��+H��晚��[��x� m�\��!�<c��T�t��=�6���b\yO��27��6��xy�xjǡPV8����LB��ѓDԺ�_\��~���^!wS�~�+�(h���q�\KJ���#;�
o����d�eF��ꍱ ����|V] j+3F�\�`�w:*�_�W�Gq�M�<�Yw���lE�_2q$�\GC��-/]�u���"�i����o��҉<zU3M��G�A;M��ޞ#}���[���5�0�t���G
4��@��@B 窋J,���DJ"����Q0c��r�TY#cJ�h�D�v�@������b��X��G��`�������/�S�;L�����o�ۍ��X�瑜�Rm܆�����V^�Qe^p�����u)�g~��׉"Wf��n
	'��M�K6�l񿆫c �N�Y8;�>��gJj%]<�=crW$^�v�@�~�䢶��1C	ι
%������yx�F������k�B�s�ޔ�?�>�����X];	,��+�yɉ���S��Z*��3]���B� i����B�f�6|�H�k���q�<H���aO*?��fO �J_��*(��s	 R�|t��Q�(��q�?	ZZw�F0?�G����?7�;�}�+zB�ms���',�膶,H�v"�/�>�ϜB���l!+��Qr��NAA٭ [�w)��9���o��9�艾K4w
�S#���/�S�s���.kp)ky>֜�gw��%�����JN!X�.�O/;)�f�/��&3wX.������&,��:��m�:�S,IeGL)����*��0|����k.h,��p��zE��Rf�l��ЌR���hp\h�Vm�&Z�D������)"�C���5pR��	欒'����ƈ�=v�㘵�!��̒��.�%������dd��sDH,��ߛ�V`��C����gA��#���g��kdA\0+����q#�6+d�e��"t��jg�Q^IT����/i��~�&>���@k(4���ϊ��u)����
WxR݉7j�K�Q�?��B�x:!��X�����2�	������װ;�0� #�/yvlգ�|!�r݁P��>�`
ٛ	o/o� iwދ0P3s��6�^�c����)��澤+�uK1u��a�
� ����#���o����7���OCQ]����>�T8n���ܻ����x�C-�s"DD;�a��Z).��<O���&Ll���֧-����sn`~&�Y����&��d�9I�13(��0���h�6�w��lG|-]��.��:�y�H���h��D����t1����߃�꒼�A���3-�w�uF��}���m���/ݽ`i"�(/�0V��)(c#{��L�h>�d�I���U�g/�;'��}S��?�J�#uTv�Ad�bss�;��2��s�A~�|]�����V��6����쀺U���s\�P��1h��o�N1�v�p�K�B�`���|�.0a�뽑���\��с9Ɋ�2���o�A�\�� m\�&�x����A�wz�N]~��=C��X.3�����Vh,ؓ�R�ї�ƀz�$<����e����0XĄ
7̚�4�z0�$T�cW[Ma��w�ץ]T���{���H�|��=�e|7�L+*�v�:�d�1����F�am ���]���)�8���&0�+k��|f�-��$��[7³Fwz�\@ͼ/�eGo��3���nzLV�fe�3�B�\1�
�x����d�В҃�R�}T���S��lͫ�I�)�����/<�Lf�ϴk=����� �4΂6A>�n<L�d�Q���C%l�οء܎2�"oڗ.뺄h}�U����ɱf困��YS-��H6ϟ
�H��-47�tz�C+J��nH����to_��;�8cs�TR-�'��<^u��)��A� �`~+��>B��z��+��Z
�߂a�})vW��Hg���27tb���3��Z�X�����0M��neb�<�'4*�f&ʛ����_��`V=s"/����1_�Շp �X�KUU½�k�<=�8�ќ^�����:?A������ā�Q蛪�q�cN"�O'	Tg�$uw����=��@Lϼ��2�=�I����M D�L��;�Sg��R?ӹ��Z�i;���V�g7>ڋ��-=���
�ڄ5p%�tA];�A��g�궦���X��M ��Y����_o�6#=�ؗɵ��ͺ�����6!Ԅ��E<NEܱk��yiA������9O�M9M�E�n��>�i�d�,���23��������ۼ��rg�rԗ�V�%{U����f�o�e��5�ZE�<�C�u�ދ�}7u"�f��a����9���F}�����Ħ(�HC��B/)�A�)�Ց��{Q�T�,	���o�E�3j�A�(��6��J��8�nD�C�����?FE�Ǫ�c(�����a�[�x� .�I���	ǈ���ڛ�b_��H�N�B�nѤ.�rȽv�\S;�	���#t�v�s��t�;zY��N��$��� J��(F�A���`�N-�V!����/|�'�[�䢄RU��9�3w�2���fD�x�Z�
��e����P��&��8���E���e!��]��y҃�$���qƅ-^7��
�XXY9�)2(�M,����gF�l��ұ�����'ַ�D�nچ�u�TH3p$�`��	��i����v��������!]��d�t~%H��T�|`�lw�5�@2/c�jl�m٧��n�a
5`�`�l�T�egR�x��3"�[Q��^��-�'�����C�r�t[�y�&��(Bl�
 ���z���{�A���l��S��]/Q�K��o)7-H�t@����J���W��r}�O�k�^=/��F^o\�"<(��g��($��{)]X*$�Q��� ޔ� pI$w+�$��\z<1���	���"f��W�PCj�5p6Ӽ����{�3J$�SŮdc�#6��P �M��kr*ϖ=�N��uQ�d��4L'��dd{\��g�{�b�������������'�0�Yɉf��׹��ۗUmJ!���)I�@��?km�S�n������;$��ۦ�����M�o{��m���?y_>�8���l�Q��x6��?jSds�ɦ���Z����Y�	�@�ۛ ������!�LV$���*`�s�K���z�Bl���߽��2Qcqe����$�+i���4 �<���s�X8c{����9�<Y�E�^-=@.��w�9��j�@ܡM�S����ī�Q�<�=A�*ݖP�~���8.�ݍlH<�(���HV�&-f�{5Gr�+vw���Zh5�6�=?���b��!g1H�Úu�0h�`$���u�)�4��@�5o�:x>���W�F���L�v y�HALvB�s����+�X�G�!�u���ςN�(��IU��OۣQ��tv���n��d[��J�o����x��!Î�I~b��UcS&P�2CBj�N2ۦ�&@�*qƐC�x��i�Gͯ=-h�q�!2h��{p�b ���H�P'�@�� �"؃:��|GGA�G��Y>/�{LZ���F��ʞx��5 &���ŧ ��QkP���B[W!H���=/������2���I�o�S6�As��k>���uG\H��(�KfNr�d�AO����,�c8�:����mT��.�vq��������΃�g�d�c�tVg=j�_
�=T����}|A�?RP2���1/4������v����1����@&�WV��V����iIl�̞Kn��E5��N�OF��B$�z�/�}�T��՗�(�c`Q}I#qS-�x~��?:2��A�n�1�a����l̳H)�N"l*Oy�zν�o�|�/�E�4m��t g�����o��	���n��<��X�JTڀ �\#y�I%<�qJHu��h_�(``�`���5���Ӛ�ܻAZOg���`���SyhrFZ���ٚ�탸�k���{�ú�3W��weE�#+[F�	���#�h�J��@�!��3(�Đ�Fz%����J�$e�������"�����$��ѿ��Xqf!/�s,j��>�gE*�fK{tn�&���1���M�#���R+uG#�V�z�X��V��$�{�N?���f��XV͙�Yi�����P�ȋ	Jx2�ۚ�=>��ײ��Tu,9�v�7d��˚x
_��q������dvxf0y�Y������Ԟ�l�j� ��`T�x^ð>0��g��_�}y�
W�PK�/�iq9m�1��������S|��0�$��$N����-D�Dan��6)V�3�[��'E����?!"��%j�f4���hw������7�l�	�#����ԭUD�qp���K}���}[	����ڎ{[s�p��i�Ɠ��~f�;Ym�Q�k��~����"Swf��?Dm����`�e˾^��LS1e�}lP;v.#f�S3���o{�iB0�B,w���7�����2���%�=���Q�n	:��9˧{�#gt��?��䁠�
K�����#���]�"����w�a��F�1�D�V\�2���](xp���>:?����rI\��u;�s��Z��OiJz6�O�v�Ecӯ*����V�־LDO+v�bX�cŗf���k�>c�8ʴ��O&����|+]`|��Z�uB�T�a� ?<�1l���xޓ�#[K֞B���H��&C!0��*�l>㱎�Z��\ǑwlD)+6N��.8�x����V�D�v��\�/�^{,*�8)`lˍ3ٴ����I�-�K� �Uz+f¡R��j�*�������/P��ġ���ɫdbSw�fǇ/��O�{0/�8f_E�Qy�-���:���\�z�Ƣ6f����'Ytl�����wF��]���H� �G]�T��Wo/�g�:H�/û`����Dh#@������K�Ŗ�K�vƾ�x�A� k�"��e)2ȗ<�kV>UyaVT�w���+gc.w���=�(̩�Ea��-�?DL�q�a��9�!{o�S^&����r��_���ş��=�"�����O�Y�rY.9� B�*����d�kM�����զ��H�3�s^&VM�D�Z�����=�򅩟	
]^�<6�����/�D&�#�Ϙ.b�Lg7�s~���,ؙ�s�D�A�-��%��bY�
^��O���,�ӮǭR
�%g-S�FOԬ���52��͹'��#������T	a���W�����= ?x�b���k����N��X��m�=/es+r[�*K�#��N��s�0kb8>>Ԍpˋ���U-�V����wo���	cD+�K	��3$�p>j�pp�of�3!�t�nV���w����Z�48��f%)�e���n��O�)�<R{4���'/�����pAe��(�yT�֨b�}��IzG��9JT?&?���9�>��Q�]٤�za?I����d�������@�*=ʁ��p��2�/r�~3K@�}���(8��'��l�!�֩�jP<��p�$4�1�2'�f�O����r��et&�~mtaS� \#��u�喂�?4�5|G�{�@�)�e��[ ��ft˾�}��ݘtI���y���F�Mϓ��b�Fg�h���o��FT!wF�p/xI��4�;�����4h5�n�HrҠe���(kϠdt��W�	�S%�n�T�w���*RT)��-��S������<����]͞^w"��L[BW�HVZ�/�ۣO�aKK��`������X�(>����o��% z����=��K�  ���Um`,��(sQ�Z=7*B��(��բ�W,�-���ǆ�|��T��,�'^/Z��r�>��)Z�|��dB�
/0��{
��}�T~[5�Ɂ5)�F�)��R�ZA�qJn^x�n|�{��D��'����8��֔(
5�IW����Gը���a��rv�1b�M��+�C����[b�Խ0�eWJWֳX�U�������
�fl�����<������`�NK��Fo"!�d~m�z�����k���X@d��F4�!=���j�b_g��H���93��]��.�(��7?�P#^���V2D�u�@p��Vx���3䍅���������B�A΋�.��X��9;]�!4wO	(.҉l��)94��|$#�5âKK���P�-�Y�g�~�o䉊JV��0�#�CzO)GdWfr�������P*k6���s9v� ��q/��6��'��c�\�_?Ȥ��]+���`
)t>w$}����y���`&��Q���oՇ2��Ԓ��D��F�`�W��O��h��чo�,�fΧv�T���̚���>Q�1�J+��xץc�TuC��+��Hbvn8��D���+�e&�,!\��7��E�Z��|�ST��!�R��}Ɲ7�������"���7����d������#�)d�e�]�}��`��;��;4��~�H1�0v:����9����n���h�,6�KYP*X ��
���X�*"xX���E:C��G���B	WYss����&�*��wL|>��Y�{�,w�eJUKG���'��'�ĭ�ʹ��{�X��(��şc�E�ޔ�g���xD�Y4U"2d�H[Vz�x���	�\^���BV��9+|�5�(E��u��ee,�����"4�F��P��g�w�O�XL#��H����WKM�B�!tB[$+X��;zSM�g
+�l�X��?)5���򪮭+�c�g��UF}��,#�|f�ײg瓧pW�ސ�͛�Zy2�9������+�ձ#��yH~�J�80=�{m�AsmMS�8]�ȅ����Vŏ�ɯ������B�y,>Z��1�ْC��)�3$�r�Ae���h�A3�6Q>�6�����S�6��\�X�u���Q�aX1k�C��xn�eA���^���A�£���0�"V#��]\p~��N�}��EEE�� t�DC�]D�f�)1�c�*��ur���-�qD5_T�V8	�:У�W�<5e���ԗ����#��C
c�釬�����$�0�r���*TX�>��'�r���O��ō��X�d���Z7\9MIh%&j3a��b��AV���М��&����H��AtH>Kgp���~S�	G���kl:�g�s-�n
vk�S�1���v��[�ŁS٧8�XզEr�,Z�&^n�r.������
��C �〆'䜫?���hp��J����4G�@�"��U�6vi�U��W��ʩͨ"���Ģ�%;��ݘb>I�v�+b 8WDz&��YTA��.ԻDrJH�RbB�4����` �mp��6lj�ac�S��3�I#9�-�h!�R&���,h�x�z6���j�B�S� z�-��LۼuH���~{�c,wSǇ�È&���=��Rp?�:m���.��އC��_��j
�W�jCjj���a2.m&u-l�]�����I�@����j��O���6Ҷ�V���u��P��`�c��o|��ϴ��a�a���mRL�#J"(_4���Ν͋4���"#)S�#ˡ,sg����A������%������}VX���5c"<�f,������'�6��&l���R�XY�:���ϣ�]˛U�o�Y�(�gJ�FH�|�R��!PBC�Yz1�!�8�������N�D�q!䩧cJ{i��\KXK���W����si�!jy̧e)%�3�.
)lޥ$8 ?#p��~"����L�ϔkI�����@(Ӡ��	Ā�Uh����)@L�j,I.�~��cu��,�=NT!��I:f��*��� ��tP�:3`�
1���?���p�v�p�cV�E�C8Š_��1�۲�������V�+/�l�%T�������'�%J�֭����7t�FF1���L��|�M$���LK6�F���ةK���'jؚ���<^�/���1cW �^�!�k�qG �6\�3�� �W0$L�ҋ����)������Q������7S	fm����Ջ�u{��
�|б�k��P?��mI�����8�%t��*c���qt8�V�&b~�O�Ǜ����v>#`�#��%�����T(�K��e�\kY\����Q[����f� ^[s���LfJ!�+1-M�u
�����I|ǰ�|����4~	O#��f>S�'�AI��r�\�Y<U�)�?�����ES�D����p�����D/n�U4���3��imhH�t�\��
t��93��Im�����E�t�_�#w��12��4�S�E�Z�*iD2��z2� +��h�+̤�x�8~�v[z?�s
�槿%k?�)nrJ����+&8��#Z�1U��_M �I��xt�bU�)��e ����I����:;W��S6��$�1I6Ѿ`V��Q�dyկ�k�G7���¿�6 V,?�#�Ql;�6��'˒���1|�L��C�Ew�Y�z��侎�r1�~6�W(H.7�ґ��y���}Y�;Cȵ*Y�
.t�M��K(*qF�iߵV�P�2�0����#�}������s�I(�#��̒�Be�`�һ+4ۯr q��M��yqǞ,����ԩ�X6'W(b��Q�hcŘ��th܇�"R3&�3p�^>����u���۴B鮴�Z��X)���NM~X]Hn]�jÛ��f�#��O�ɢ�
�O>�4L��7ʾ�+V���3�3U8�k &�m���Q�l.�tA�j�aU�?\g�c�R�S�^�J� [ѳT[}�;;|z�~4�7/�f���\���x=�Z�-8�m���Ǎe����{�	�#��ӵ��EO}u��G���u�YB��ص�
1��<�b ;��b4��AߔV�(�=Ҋ���{��f��5(\�j%�ac�� �;��o�0)�>��.0��cM�r,=�C��$ͣ�o-�}Z�N��d�Zpx,���2k���S�dbA��تc�D�٘�/����ɞ/�����3��ٞ_Y(50�ͭ�%��v��,$�g�2�H��� ?�����l'��tۘ�d[��f�>i=9�e�^E��Jn�ݷ?���7��qK�8.	 ~w�Pf�z���{�nmPC�p�O(�{��6�1m w���n�h�K�6�CRT�P��۲)������,�utH�}��oƥ����H�b	5���'���}��U�QW(�U�$�44��y�۰j
�G&�3��[T< .�MW�Or=GNA\�z�4*I�F��Xfv9����:�����|�'�зaQ�s)K��w>���������&���jMK :����5���|����T;F�����[;�^1\v7܇��ɸB�"e�Yi�dj}2�3p���}�4�;K��CƒF�e?���@�e�
B�y��=J(Z&YGm��NzX��ԝ�D���.�9����F$�% o�Ü]��c��PF�:�.^҄�����"ྜྷub�jJ���"(�r�m!���h�Zu�~���o�T���@Uj�o26n�}����<��}��@�~S��8
�q▎�#H�x8���5��D$�q<���G�/��L����}���XPqO�5��ߎi,+����d���W�n��*5��Y�  ���j�׶^wG�P����.?V��,���P�TL;��zI	�O�e�0	��mL�7�y�s��(&I���&`��N�2xbM���F�I[f:j�o������&�.����,�g}I����@�k췸��"�c����]�3�!!ݐp	�`�h-��+���%Զ���s���h�r������#b�0a�=	��'�#"���DU��S��5]TD!�0T��e*�#F�)���(�oP�Ol��9��5�[�YD���]!��\$f�<�< ��)���^7=��l/P{{�# ���Nk'�}��9E��s�J��JOS ��Q�qc�f'PV�b#�g���v^$Jv�W�������u�[�^�R�m�u�Ygr��4=n���e4s��b�_J�M�ޢ?��V���Y�|$���Ϧ]#��Yܘ<��}�ʽi�ܳ�_co�[�k0W�5����	�"/����+�AE�(�L%�.4!Z ������=�O�C��]��Ŭ~�]�� PC�����{�L�JB���N��'�H�e+s�Ι#�=�Ϛ�T%eC覱`����H�5�e�"i	"�{s�����-�@ΰy1,L^��VoQ15������`�KX���%B�Aĉ�3�SUH�U���|f�s
pN�'K�w���ͽLЭ[ �����"$W���7r���;���������*�l-LG�q��L͠�U]�0Ai\���Fм0w%�7	 U������9%�� ����$�\e��2D6e�sn�P7���[S�G%��ڌ.u7��HuDf]#���|_�wd�Ƅ��L���I��!�D�p#�f�ېt\FEZrl_�7q���O���{�,�^h�*�=�8��LЙ��Z��� �q�uWb$M|k��6�f��� <�6�����1�e/ X@6�&BLM��I��\~ir�o���kKg��e���v ���� �D*����m �h������_h.%����M����*�!ח�7��ȡ�*7(������(@�~��V�M�}�����=�����%�x���nMuŝ�n�བྷ<���[��n��e����^)H����S�]�]�y5�G�^b=Y�1�t������9�u�mȇ6���f�߆@��ŋ~�lpA��jڽv��N=V}4��Kx���)��Ež��j]93�֚����)-F.��H�)&_D�7-��D8V�|ؿ�"iTB����ko�����u2y՞�~8r�����CrS�T����4#n�/ j׼��I������LH\��č��[������Վ���x?��ʟU�;M�Wԣi�{̗\�Z:�l#�tD7h<	�t5�Hv������r|m9���ZJǉ���W�P����}3�MQ�J���_1��ǰ9��f.�"�A9����}x�{J����e����|�K?5�K�~�^	�A�ҥ�,&74�&}�5$�Զ��I��<�u
��e*�RU��d��A8E���튐�v����3���ѫN���aS����$}7g.�؀��FuߊB#��ͭX�qۡ^��&lD�}��hSK�9i�vމl���4J�/�j�8W����U��G����K�;��~x�lt��XF*���d�jݴ@�B�U�&!`�x�ٽ����<(e��դ�.�y�����/�e��@ӛ�����������l���3@r�=��RD�`�嫩�.M�D���H�rS�T��P�÷�;��h?��?�8�s�q��@��^�!�T�"&�fL/��h�����@\HR�yS��H#	�A���g�2.�7Q���:i��ş��;u�6��A�(���㷝�$�7Y/�8��<��\��_ķ�ܓ@c���$�4Iı����g�G(9����e�A�����̪����ʙUr����ho&��T�u�s}o�&�M�&��xZ���R��\K�Q4�Ѱpz�J�:�'��[�s��o͙��P.9D��/���g��pA��k��ǜE�C�����5���2�͢��MT;���V%k�9�Qc���i�sR%��U!1 5��=g�ώ��VgC|��x��	/'E@���i"?;�<��] ڭ�\0f�rI�*���f�0B�v� V�)1p�d�'H�	���خ�JT�)YrTմ��c3l�l�ݳ����L\A�y��q�Kt��~��L�*��gWsl�%5bw�?��(P7.�)H��Z\�{�GG����l��yj� ��i�շ�-�P�"��
��	}?��Ϧ4pK/�s��p~iQ��
��7�Dg��G���� 1dW�/�>�*�׽�p��ن�N��:U����F������ @3�Mm��Z,�@jn�1o(�(z�q2���ZG�F�3KO!�B���[��ڗqo�G0[�"V�:�.01HF�Z~���˟+v�E^�EQ"����� ��2��I7̆���HRO�!���g�"�!0�v��6��@Ab#Aqv{I�7��w��&J��S��;H
�p�<��,�
c��"q�K���_x`�Hg�d��۽��->7@�d*�_f_F���Fu��-�� no�q�����Sp��݀��.r,�Ξ�P|�2�:�\G0&����fK�����.O}��c>��#���j}��W��^�HB;x��6@��r���rp6l���: H�ll�3�c���f��Y��
?Y����j�ףT4��}l@��*�z����x)���־R>5y
Ae�Z��ǓŨ:��nR��`1�p�*̟/¹���g�<�\���u��k.�%_����\��3���FU�@��Ȓ��+#�k����}��4�cu c�z*z��~��1����rL�<�Y�:�:
-�h�/u�1Μ0CA���'���d^9�
����c��z�Ut���_���U�F-�^;�)�j`�f�xa[�W����^e�w�1�C�1�T��_S����^�c-'(�,�mI�Qc��aS%L�R=pgp����j�#\���2�.��\v"�v�հ Y�����P?Y��S@Ee�㔺��@VN��^Lh'��x��z0�1��Ut�y5���/�BvģTkwuĞ�士O��;2D{���S���,�c�!������߆o�x0@���uw��%�I�/3��uT��c��7	�m-�`�/6_������>I���� �S�pBʨ?!�G�6onǹ��r�Rd��B�sK�g]-�̔n���y-���D���	#CU�-~�I�cA���I@�4l�y�Mw&��PnH�_)�D��U+<b&��[�3�ٕ~K?�Ay%SѹǊO Rd嗈m��(����r�V@�<7Y�;ԡ�k�8��N�M[�n��!��ep��uo9>���F����gT�����$���8��[���D���Y-�+�a��S��<�qi��=��n�v�[�\����Fd��y�,T,�9w�6��ԢUM|G����t���/:ND+��:�Da�Z6_8���k�(d:TX��mS]r�[g*��f�P� �pG�r1�z�9�Z�k�D��� ˪��\�K�!�&V��b�֍����l0��]9�U�80FC&�&S��I�]j�*�����1pa@"�V�X{��g��"�n��i�������O��om!T{����n������`؂Kr�� WD�]�����d�1ыt2��W�� ��F�*���#�c�rR��	� hj���1����`�Z�Ź�Jx~ka�$
 ���Ʉ*}��b��f
���TwC	���ï��`�Ȕ��Ԗ�W�d��W@op?����d��oE7�"����=���V�,,����=���Ё�w(�H�v�b����<
P��Xl���J }��E���w$����0�{� �oPމ<�D�Od��"�)ُ7�����_�3-�1�qѲ�D�L2�Z��^L0��U���l�H��_~��j��Lxp��w��2v�=z��}r��1_�BZ�w����p��v�*���LS�F�����'��+�f|�h�{K�*���+���,>,��"��qN��+^Ŷ8�.��Hn��*�o8�(��IY��p�e�^ȝ�ᵓ�[���è���X6'(PQ���կu?�����O��E!"�ћ�����m�=2�1�m�-:�h9�~���O��!L�3����֤8ʳ����I#Gǘ�wW�Ub��n�{�P+i�Xn��M����R��׽��ix�L��e�'cJ���KV�	m@���hyC��n���T`�2����Z�X�:�4%�`��FXAWB���A�u���6Ge��D���,}�cd��+���Hp�N��=aj�5`�P��Ow��<��G;�uܑu��OOn��[2�K�v��%n��r�l)e�02<�Vf�IJ��&ȋH���
�P=/��5D�T��rZ@�����U�D�d5��y>6&P��9
�������\8!<a�ݩL�����z$A��6w���@z4�z�����Y���|�X+�[x�~b(
N;���˩��M��5$c������y���B&�*��a��C)K�=�S��-F�/��3�y�v�D���H
�����W����D\=FJ�}b�91Kۃ#��ʙ���W�֟��!y�%�k��I�T#���I+�����NU�""�
����MA/]SL:`�X�E:���%Ff�Q�Ǯ*qo��l�й����'搅��)!^��k���F;�0�����NH������Rf��o�x?�[�1�DE1���=��E�"r�H!���+SV�� h_3�����	�����A��ޞ�j|-9��3G��gs	��<��gL$�wS:���u(�+����B�:f�j#`��B���w�@;#m�?H�n����w��Ȼ{w��9�2����T��6�&��m�F8r�B[�W��ýlN��� �̄r�F�r^�c]���{nB(�M����"����X� -eP{Z�0��O%L4|�c�^��}���U����T����oL)��"�{�h2K�e����.��Ǖ�~��;�jJ����?�����X~D����e;�pׅ ��������tih��$Ȑ�-��X��U�J��&S�f��� ���вX�p#�C����=�3�H`ϫj=���@���%Y�����V��:ތ�_1�_����u7̛_!�����l*�^��N�N��I���6�S�h����u�6�b(����U�*�z����q���p�s@�8tJS��G(~S*H�+�<
5�[� h�HN���@y�cd��~�}5ѝ�������TM��~��*�%�]~��y�(,�cU�_���e���i=�T>�T���ҸG-F�!�$� VU��S(���O�}(�|G�}�ci�O5h����!�nH �gƘ9.!��sx.�
5�Hy��0�(�6[0S���2MﭙT��E_��I\x��I�]&��<�U^F�p�Z�h)�}[�R}�/�xQ{�� ������o�����{m^��/�də_=+D�i�b̔�W�`d��eA@��t�t��Z�yɆ-�RxF�&�]Q����3���/��&P�ƈ+����Ϙ��=Ch�5���6�U�)��k���\KZ~�P��Y�y�� ~��k.�yL}���$\�G8�R,�#o��[�c�*̄k]$�t�e	c¼�<!�G��nf����L28�]?7���Q� ܂ ]Z��B�y��r� ���n��~ �R����}��	c���S�*��R
d�ѿҞajw��q�!A7±�4%����	KA��i-��2V�Fj㗠�t �nXj4�0�RŖqz�g��Iw�F
B����k���e>��nW�Xr_�*w�3|*��Zs.�y:<Gb��e�<Jxp����寛뢬3����^���e�V?n��.Y�Fl����统�f�]-=�ng٘���]���ÂQ9����EP.�Xd��ڈ�/�5XϷ3�Drt�"�.i
qJ��ƕ��3�J@�2OHpo,�v��'v�(K�#yL�iX�f(�o��U��^����0��v8�1y�w���A�y!�e�|+��(o�rk��nsgSc��~NJ��p�d�Wo�Xؙc4f�Ԕ�WF�v����#n���|��4C#��*f+����~?ɀ���S��*V35�����bb��a�s�xS�M�S��I����ޱ+,��Y�}	��%Z�X������}�9�6N��"��~Da�3z�Lh��[I�qw}hLh��.�R�$ڀ���咙$`5�SJ�Ykt섗�S�g���>���q$����x���q���	����vcGj��$�-���[I�O2�F(U@�6K��܂�b�c|��C��쑾� �{�8���*���!E�����6�Ȫi1����-�8\�1s⧞9��ߠ�����G��*09&�v�#�X1��6;�@~_Qv�!�@��6�{�V��۶�Wp���[z��@48u��L�nu��-��X�{Ԋv�eg���;vk5������-�Jvtn�&�lV�6��<M��%��+����rה���bl:B�6Z�� K�NcLQ���tC��s➛���y�t�ߺ��'����,#�{8Ng�'��v�r>ULpْM"��*=�6��Zd�8��-�
Q��T��{.�ď���G-�):yp���j��[�QCjUs�V#� ����T�0�J�;�YZ�>��f��Xz/Gk2c]���=�H��(�F11��AM�.{B� �m#�y�2��/���������7���&� �t,��? 5MIX�C�	t�� ��]d4�!�T]B8��� �áƢ{�ȁx����f%���>({a�wp��B�;�+�%ON�Uʉ���%���.iu�
q��L�9���lb�:/�0�ě`'�X<��b�P�m��[��aQʹ&�nv%�߃5�F��NF�K����?�_�FߌC݉��v��8����|�*�[,H2��K1s8u�c�Tڕ�io�-i)����ѱ�,�NZ����B^m2_m���⚙�ąPG��x>�����C�縂K7&D��sq8���]����K<����2���إ}¨�R@�ݼ��}�'V�8!?��]3��,�j}jpl���-k�c�9��W/:y)�5�Z���8�����j��Q�DIY=ԉ��e]�="�k�_m�DuJ����� ��Sd�}�R+��)Y�5>~�An���\�j]��ZI����\T��~-	��O�z��J13��= r	$P��P�@ƌ���NJ|}��]�T�뿧�m8�h�5���E�U�j�\��;"1��#r��I�:�dO�u��NQ�D� �o�D�E��Aџǜ���[��J0j�f0���lX�$X��`D|°��P�{z[�l��H;��� ��0A2O�DZ�˾��P�v��G���vH�9[�o�;������L6���fG����0��_�Z�8�#Qj߀�V��Ț�����%?�����Q*ؤʎW�DNUa�4gb	�$,s�U�69E[w�}��ъw+(eh�}z/����;Kl�2[���]�UNO%��K�Fbz��)�F~۸�(�W�=�m�*8�yCs�(��7D��M����ùf�-�A��h�PF3'�N����.���A���K2�I���=����4����@���
����~�A9�#?�F�?��#!4�������ti�!8JW���	����^u���t���:�����D(�iM����Q1 s�%Z��L�@�j.�Qk��1�u@'���C�&�u�;9O�I\�ր��+4��6ţ��"�4hK@��v�͘����T?r/�������-1��pK��0/}H��:��O�2���(ͫ�7�J�F�a�*gi=��B�`���0r�#*z�!�fK��	��3��B�u�� �1��ؤ8M6��������Ẋ�Q�E+b��E����L�F�b�J�e$�����2�f�I�O���WVNlj�����m���	���(��N�	�����F�V~[=�T���B���ӎU�n~V;���}����9a�k�d��+C��ml30R�j
B��1,6أ���|�u�����v@�B�i��W������:����+Az��=�qRd��I�+����)�M�h�]�
.���R�D�%1MĀCSp�Ύ}Z,Ec��+�:s���%Ւ,*/ɜF��p?G䟦�O�2�K���M���W�C�k�j�u[B�a�iظ�����A>:��n����>��Q�ȍ���p/�0�mu��1�*z+D\�ͅ��Y�%�L����T�[�������W\��ZB!�
 *�Y��A�N�%%{�T������)���4�����'�o��V��WB��.?u���~<:RV��(7�{!t+C�?v��BM�?K"��t+�8k
���b&)��q�i��+���������Q��Ȣ����,dr-?�hޮ�է�,��d6�Tj$��a���ˉ��9�-m��.8�}�ր�6��Ez�K4�r	�?����-�d�ߗ�\9fA�`Ѓ��ߖ!g,D��UO�q!�8֞]��2Ծ�&��Cx�{�T�,s��˕ X�dP��6�����~��W�I�IUZ��>P?���G�f�yk�c�um�0N�:�������-�Q#:�ymZ{)(�
�yh�7ø������1��n6���E.�ܵ�8,���<6����7�����G����˲wlL��k�^�w��<�?%�G3�e����%mq���Y�;��'��2嵉K*m���yV�
M�Oa|�9�\�DD�my�a��Se�R��T�J��
�r��p�G���:�.�� ]�)im[����j��2%th�7{AA���>�;�o�ހ�����h�^Ϯe�Mlʉ�r!���l���KWs$��tj��^���$�JgwXqH�%�����QC)��ZI�(N����x?�:�4)Q�c�����oK����erC��k�F��S���_�"��.�Q1�'�Jyn�"�#/h��9cYS�2�t�A���+��&�*��M�\�OB���w��.��M�筢�RH��P.�g�������LNtם�z9>��`���ܑv����笯����)�-��ʇ�m
DI�&t�����t���u�|6r�\������Ȉ���T�>j�H�֛^���[��o���XI�zRH�r�iit��Y5��X��l~��6ƙWU/h�{n�4WLԮdh1���8Z�O [���� qU�íb�ng���ı��4���H�q�}@�h0]l��BL���T�i�є%����U D�/"��jO.��Ȳ�#��K.�Ho�*h��6 
㗕��R��t�"��0���۠��]9�'�;�\�4�~�'���(˅*Y��V�O�T��|C��L?�AV=��a�>˅I2"ߒy�Bʷ��4��U��a��M�ɈJ����\��Y SE���E#Fh2>�N��"��rWܞ~��tŵ�&�d�����[��˾Y�wok�j�AI�jR����>q��r�3<��C�ѩ���Ի'��Ғ�%�s,m��Μ�{�*ܣ	sNfK����T�jc(���#���ů��>���`]����p���&�#Ð�����8����K��Uc������nD�o;ŉ ����pc��-*kT4�Ry���]�4�h��KB(�R�h�N�C�F�]0*Z��Ugq ��N�&8��z�l.eK}�	%O�5b%P $!{���N�Q��Q?^�F�E���+q+��]� G�r��jNq�0������T��6�u �޿�k�[z��컉�#��'v�h�<x�髛I8�ZC���⎯"�a���b�nVV��pZ�Ƌ?�5�9���j��_J3�1ӱ��Q�Q���;�L�]����|��3��ʰ�3����C��������f�)P`�8�+�l-k�?�!;�k~5�4�҂��v�W�qe�Nq.�i7&`'��2�<�y��iZz���PQz��|�p�:d�*W�zr~x\��YG����w�ob
�c��H���;48r�
�q&k�̎)���sH�\�z�qOޅ��^m��e���E��0�s#Ax _����^9>��v����ȕ;J:���?�X69|�����P�])N����L�����/޲x�@񜉁χFQT�d�m�_d�W95�D	p�1���P�Y�X~8�������1�O���=�'��`�"
����Xն��#�ފ���&��0�/��O~id�$j׽��*��l�t���n�BF	��v�|��Ǐ]��)�wS)	?��US��)�HH�o��*�Y�ؼ���N��؝��q��ǍӓmX��爾+ȪhL�K��sY��j� ��f��KJ�|VL�Ag� �;��G<��@j���E��������'�tǩ����K�j�Eѡ�����cZ�$���X��f�4��^��l��#�*�U�:�N�/V'�aڱ�F� ��Bn�9k6�5����.N�-R�0
F�o�8E����6y�޼�=�J,چ��{zb������������.����1V�7<�7�1*�����VL��¬Љ-9"�� ���kȗ�IG�֏�"�|����I��e���ꐪ��:;��amU�d]����C./�hQL�e�_G���q��q�;N�S�������ʮ;��V���C�շ��Y�l�4�e���oyNl��V[�g��4߰�^E��ߝ�Gw�L$gxM���2���~r��h�J~g��5>�:���=�2)#�("ܘ���Mv�t$�X�LUa�G��%5x3�w�q������]���Kh�ITG}A���u��P�v�&;�Cu��1�"zsÀ��>:�s���9��Ed�Ӷ�K��Tu[�永���7C��`L�����ȱ��w����(r��>8�CT���V¹@_U��aд�~VH�2�U��`�`]��[��+5�Y3)a�@���*�3��	LE�I|����B��^�juay��������!A@��j����p'�`�d��vCi}F&��cA�k�|M�Q�e8��8qJ��t�-`c3ߘ�L�L;�t��M�� |�Ȯ�J���3uS�AIp��P�զ0���m�O����\�����!�H�eL��jG�)�_QP�}~F�M��F9]3��f������r2��L}H| Ł��Y9�ڇ��[�~c\�
wgl��ԉ�U%�c��V+��<l���`��5�����1x��!��֣ݼuU
���}5ݧ�:�]06������j��U¨��[�۬L�Δt�j3w�a(4�(<��I�H�����IA���F�B�/xEs�﨎	i����a���HӜCq�j�����[^Ƃd �n����>�}�LiE��)C�������@��`{�܂,�L�{�!T��/����k����3 ^;h�J`��� 2�^!��~}��5-�8��]|dP�TۖP UZa�1���t���o��'�H:�`���,�#BJ�Al$��<p���j�,�#;8d,#Rv	fδ"�$�m���]~P���:ѳZ�^��^7��W_�{mů�.�&ٽ-��QD���C9�f"�ꍞ%����J����io29�A��-]q�&z���>���U/n�2��)F�)��NCAc�D���JAP=];C��ᦳ+�>d���oa��&N���P���[����^���Q��zd*P�ߟ�&�H�C���z��3�<��xc�@�+�S��cEte3���������Iňؐv��q����7�}D�؟�X��|��=�r���]�l���͚�-��t��o�y+$9���k�}޾�<�G	��BBP�Ev{���h_��E!�q��������g���*�/��Jx�ʍ�`�bK�?��5=cu`�@̓�������S�(�{m���dhz���Sx)sr��ٝ��/4�b�p3YκT�ec��M�¡06B҄�=7QTThI�T ��j��������p̈́bfm�\	���(f���C�-����� ����T+wywg���������cc�}�`z��b$w!{)٪�$�;cKQ/c2#�1��1[�%;�/�f���h42
�kd@��8=���6��p�qi�7�N�o{��~][p]RN{�YͫY"���Z��y�wh�{��q_�S7#0s�w4P@�+S��+����m�Z���V�ݻ!�����Ӗ6l�>�����qX�`v���S9M0�֨��|�Uq{��.{�n�a�e#�^A% ���B����I-����s�I�Z�'H�L#�T�F�k4(��\���/]�R3i.�R�`��	��J�(l�Y3��b����(I)������q��ۮ������C��� u/��T&�7У:��F�?��|*I��ꡭ�*��/Q�hG��UhAZ�ք<]�fe��vH~��f��<�������@�C�8���W���"�� ���S�a����d�0�����$ǵS��>�U�D�2A������_�P��k�.��>�h��v�([���ޕaR��a��XX�g�
��A�!�"��H��R��P���ס*3pc�C8�Ϙ���YX��s4�*$0�Qսu��S#J�V��d��s�~1�O��2�%04�+�}o�\�E�o]��/D�h��v���ʱ �>X�o�EKMz�h��"�t{���u�g���-���8�����������q��]�Y?�*f�. �+��>K�q*�t���Ag0
�fdj,A�Y�˨E�[G����&��v��b�L�G�>v� ����ǰb�[@~��4y�Z<��R]��>��ww3����'��؇����֝�9��kM��Lb�X�
�0�Ә�}&��Ay����J+��qJ��#��~���j\D{���J}���Q�1���}e /�-�+��P����;AoA�a|�vh�9欨�s1qJo3&=<`�<!>���0�����l'��k>�2��x��@���8WH1�:&-�
��FP����˕��4���čw�	��������J��Ȁ=���B&�2�Z�����c/��˺��]���і7�YTE,��%�1���ML;ئI#S�3��9�ڣ����|��و(|f�5�W �t�(��>$�u�#�:�ۣͿ6�d�pD��Z��F�����Oа�Hq�Nfhp�j��s��<��@�����wi�9C�m��^�Њ�}�%�+U���i$�X#y_�� (Z�xߘ콐Ñ�[}����g��A�V�Z��=7��� gN�����r�s�AV>g@y^jL2�o��#��E��<�'R��@t��vgh2#�ٌ�[1���Z��
�!��7s������>�p��F���L��H���|	��[Ǆ{�����G�l��@Z�Y��;y�R<a�b�.�׻x$<By\zW�ۅ�zCO���7��A���E@&�z�7&�蓯$�0�[�. Q@_�L�
�q��(�H��v��g�kR�4�0�߬�0���T_����f�L��<��S��Ph ��tk�h���?�JΖ��B� ����x&*������;R��zy{��$��L��/�h���s������fo�>�d7���nE䵴�<�O}x8qN��}dL����߫M��U6�����X�g4G�5G}��a^��t�@L%.���Q�W��/T�~��MY�$S	��������M�R�;��Cf���Шio�B�O�$�b������DR��x'g��S�p����^�'-E�^U�o�h��:���b�r(ҥ��=���U�֩�ϓ�T��T_T~1�A,�ji��S� ��̯��ޑ{�*�ڹ���y�\��6�"g���Vl�����f�n��hg���*j��ʡ���#L��^ �H�fw~yۃ�RP�4ؒ���h�$2=�����o<C�P�^���WV��w)D���~�11p�;�J$��J"9��g�1�P���;��[��ͨ���s՜�M>x����P� �캑��\ʽ����A��!�&�]<�Q�nY#�6���^�������
FF������k1Ƃ�L�%�ю�V�x�;Ƕg?�7XU'�3<����mI�Ϣ_.�so�Ld�.�{����*��]�68*p��3(�R�J|��
ij���q��q�u�q7��y�Y�d���v�H��#��4b� !��ǔZ�^D��8{�����K%�v��*S"�x��&�%z/� �~�g��Lyaw~̗��Y'zȓ�3�|�j�K��$yZa6���rF@��>��'u�+�~����K���sq���0.�ORSg�m���[��a�02���$�:Sz���V�	���1�k���SFm�Ia� ���ƙd��o�'?�� �o�%3nk�Z���O�wT}���q�|��ܿ���l��#u'���У�Y)vB��f�Q"�t���	ӫ=�X���4�ݨd)e�e�ɞ�e�Y�S��Qݹ�1A�҈Zᐬ��,ՀY+T���B%[�����������Ť��{U�n�D��� �{�Z%W6���GӼ��ƞ}�DC����ج �p�<*�n7�zҭ܍7AO��0�5͠B�x�����cGƹ8U�b�*�Qe���:_}MIW��#�wq{-�Z� (c��__GF���y5�Ct���)Nt;���
e��y�䖐ᑺ��89t����y��������+��t��%mv5��Gض6�&�(���}YD���"t�Q�C~"�)��Ԋ���5z\[iR�ρ�0�6 �f����YT�e_���-�z�iQ���tu[Ʈru{8￤S�h`])�����E��Y���iX+gTqi�x�Ù���z\�����k�S�y
`�bUϓ���DsS���}��m5����Y�l�~��b�wF����d���^�rA�K�J������ s��7�=����(!?bOo��G��n9>Z�+��ƌ~kƃ,	s0�gX���(�����(�h0��͏�����s��v6.Jnĵm��_h9Lk(ܘ��|6	|��5p�1�->r�T��*,=�mK��h#� 8r����Y`9R����m�*������?=K]���,��@fZ��_�E���?���q�S���ʎqvo���d��b���6 �E,%�=�Ӂϔ����vd�lym@�+�Jq5;��K�=��۠4wU7��䠱��W���rm�W�IP�mV���F�Qrk�"Q���䛂�v���Kl$-~<�LW�L�Y[Ƴ���`)��\�X���[N�jb����m��R��n���>"�'gr�c�8����UbG^N��4�3Cש���Zc�".�.�\��!zm~�h�kC��d�*��?g�%A۱&����r�3�T�∲-��z�M0M�P�:y�� נϴ��i�hJNq"K�$l��,H@تcY���t G"KZܠ�2UuQw?�(��Ǭ�{\�ɭ� �4G����3I�W ��Ru��83���l-����H|����/y1�[�+#�+b�!�P�%�II��� 6�J�1���"��fR*�c�=��%UHBv�xC־G;0X���S��������ĉ=������v����P^0�:ʶm�����0�z+��"a@_x}6�,���FƋ���h��YL�˻��/�:��c�|x��"c�ߚ�Yķ}��v��X�,��\)2#�G�'�<��S,]0�g�D&ttL��âXU��2���ı&��k-E<�
nHZy����|�J� h����O�_�|�ì�A�Q9�[o &��"���H|..��Pm��Br�4i1�U�#�M�@��$�.q����N��8�ωȉ.*�J%Z�� ~8h�/������`�Λ򨆻S̚�m�q�_���#��h2��1���*�8�_K~�_a��Jk!	���m��*d,#���F� �S��#l�46m��52��	��^#���ѱ����%汀�M�1(�p���l�5g>w�VkP��{i�jR؋����ϱy�#���3��������n��n�l}~Wb��N9��^�����JT�L�R��@�7��A*�� ���N�fC�*'��P��� �r�:Z���*��҃�v��s�YE �g�c§Ә;�N��CA<����=w��%��b�p������T�u���"�F|.�l-�i�62	�xʜ��,��#��a�7Pb�<���ZVj`�V���8xzҢ���M�O�����(�O�ˮ��\Ld�O�h(an.��,nW!�1ݕ6��e߹��!W^`�0�ξ;��q6���l	�� I����dK�ub���@��Ȥ*�CIP|8�o1j�3J, R�	��~�H��u�����uߝx=��9����Ga������_G�*l��Ԃ���%'��Z�ǟM�a�`n��$��z�Բ9ʓN��97�z\�H±��ѫoi!c?���U��<�ş����`�o��;v�7�H��:([>[~�}]�{��S�`�Ž�)���v�P�Q.���� -`V���Tm�hi\q8*�^I���grP�{J3A��O�UT��ŉUݾ`�6������#QГp�y31벋���yx݌ϫ��R��߃��M���_�O_�yJZ2�ߎ��F�Gz�Ȇ'{�v���㧏�u�Z���*�|
�PUXO-?�V(4BuqZW���|*,������i�s�)у�m�3q��/�ڨA��'��?���� �F3i��q��L�Ӎ��b���),���=�B�?h"��D����M�>Uo�����f"��ߌ� �����x�+�AB��=�9���B��.�t5㲠�jF-W�=[�,�Ç:d�߮R�����E�N�V�ӆI��7i&y�I��aH�"�8����8����D�_�Q�N8S�}��~�a|��C	�ݫ�hAr���7y��2�[}W濳%/$��V���,Eqgi��	�����V���L��Iu��|�F<�ٔ�;�@*˳\ȷ���p���YgN��?���w̐>�����(	/��5����N�ʱҦ�^�p�A�LWej�ܧ�+a��WݱzC`3`�'
B�,_<�[��CZ���k*O-�|�ھpWIކ��:����ZkL+(���	�4s08�w�S���>�\n�R���wK���k��Z�RT�&&�Ѩ9EM<��i�3�;}���p %;tNh�%�@ƬP����1��Rlq��򊝮O|]�}��wS���	��F ҫ|�͑�Ü6��7f����MG�Z^��no�vx�|��v�$���I� ���M��X�����ME�9~b3��\ �0������Q�~�n�x����*Au��zb�6�De��?;͹e>���˥5�$�OS�NX�\��?)n��j�nG]s�-n�oG�X���`�4�C=�����7�K)�����<�9�c�y��-NY�Ё���GnZ��ti���Q��}�s�Y�,miև��p�H~=�����tE��
L��{G����>ϴ�������k+�B�۠�N�]��L9���|�GN�ʼ���[ �m���ik��Rm��e8h  �4Z��w��1p��c�\�eoi<���\��m9&pP��y� ��D��M�C�S�qbwp�zl�;���:�6�*�y~�y�K�ȜL1H�	H2��؛,��hK5	�����2\|��t91Ge��edۦ����6��WE��n#>Y�c�XތMZ��#]�TplCr��&�{����7+�+;�0��!��Mw�w�L�&G@�p�W Qи�j����.A�)�U�hZ�_�}oǈ�YӨ�����zi�6�����+c�I��h~#���%����(�b�u"�m���u��H�҇d+�9*>����]�Y���I�-�k>�3���?|�ȂX� �O!��w����ޠ��]�ԺRxs���� Ԣ<�+��EQ |U�H	��$
����:v��6̪��y	��(�W���0�?��{�D����I8L���R+�I����fʵb�8���e`���=g�)�_�k��j� �}�A5G?3K�r�	�E&:�%vZ�L>nL�n����n.��Ę%��g���;-��F����)w}���pi@�����ČKByK�~jN:��8��n�m7
�:e�H��v\œ��.r\�;�B�����4�l���%��{H� 	 ��t�Y�����eUe'�b���|ug>ν(�[��w{
�	�.z-�4��3䩀/"���3�j����ܥ.c+g�ME�e+���h%�([�Q�iE�?(M��i����}�{�`}��M���Tt�>�Op�6]-��6�����{X8L-1�0�t�hO��p%���t�L~�X�J��E{�!�{ZDE��0�T�W�~��Q�'>8�a1��i�J�_Oa��v>�]-�(�ʓM|4L�Tb�ElL(�6��eg�\fOn��i�,��'�i����J��U�z���DvC��f�h�a!���|��y.3`�����{��V�b��g��+s�/�m���U��}hk��O%���LR�̬������:K.+	�����%��J ��`�2d�p�Ⱥpy�P�u�������������.(A�0������*�V����F:o�UC�3��ֿ
�FQ��[��9�z1¾�&�%7 �w ��<G�[]"l�x�#��Q����mp^��.\���V`���ǅU-hB�����������ĉ��\�d�?/pw�IܮZW�$�^��X�K�X*���R'��	j0K�, 6,5�#�)0���BB퀟��Cw���e�T?������)nP�����Xz�(ӣ�Eӈ�]�7G�&A�$����"�u��wo�䵸s z/�9}	�s�jma�p��/xB��'.>IO��J99s�B�ɺ�1�u!�5J�n�}t>��0!�X92l�\�� �ڤX�6��P p?�6�Q���μn�.�F5����<���4�Zf����d��7L�a#Cԣ�D��J�]���Or��n΀5�'��o�m�9�&���>�H�@B�fQ(0�"�X?UJ���wo��d\M��ߊ��h�vsz���|'S�)ۙ���$��SRq���YU�W�(V��a�M6���Y����Hs�v�Z��-Aޣ/��&N*��j(���̻��D��V�]��(=Uq>����J7w�&/DL�.�����l_�d�yюkx����E�����P���|�IRk�L�����_n}5�P/\�`}��h^ ��Z ��׊#s;N�&�M��Nц���a�7�	�`O�	�'deDٽ�D�f>w1��k��X���s�S�r�1�-`-�t�:)��Q�F�'�l7�x�A�z�����I����"�Ʉ������V&�T��[�>`�_��V�<tF���p�]W�`�]��
3�@��#�2�.Ӝ�WI��g�B�F�!�	$d����qd����s"e4�o�ӑ���Z�}J����Ixۿ߫:J0�(8o�67�b`4�^&��}�Q��d�!�4�C��B�y��y�ޠM-M4���J=��_!��(���sL�\`t�� �	zB�}�g�mg%�1�����7���I�纊��Oҳ@�Boe=��1������#/*�LZ&��}ơh�������ЏR	��K��k�)4>J�uCMqM0;�gk��}ĪK���k͐����i��#Pjt,��#j�韟�]um7|xKIlQI=����=-"�������k�S]b�<��� 4e��?�� m����cMeooj���S�>�)�#>)�J��*H݀�</��wk5�f'\���Jl�NJ�w�t�n�Ű���j^����Y~NV��<ݗ+��-�Ru�@CH���%��"�߸�����c��<�s���n5�Bم$y�L Y���_QAUy
����bn�Y'}������˷��W�H��l*�u�{�9 S�S���	�c�˪RJ��Ό��R侊z��uv(�i`�>����\�b�s�E�&;?�Wv���!�2�ّ*��Ks����
��\D������2��瀳�m�]�$]�2��v���6]}�w�a��f��^4�  n�s�W{�D<��/*؀׿�:���KA_�"yQ�����;(F���4�c�}�;�=��bꓱ�����iHS����sj`*F���C�Q��	���䘹���>u�	�kk&��A��A�+A�)���\�U ��>#���0��N;�8j�m{a�\�[��@~�l�	5���%3*⬁ʭ��&��Q;����]a�wIx�V(���vW"�>�����vwꎸ���'X�g�@����0���Phv�0L^�=[�T i`��ٶ����u��N�N�,���OyW�#��U8Q��5��}֥���Xk�Z��2C-�&Ylw�`6L�x�eO����	�*7�|=7�e:9�hF�!;��b�o�0qa�\M��l���Xjj��$u�&��wzZ� ��L�_=��xXVxJ>z6��<�(�vty��<�i�� =��tz�ɣ@5ppX�8�1��8���l���`���4��U �i=���2Җ�Xe�SQ�Ԣ��B~h���e����$X�֒
ݑT��p��O��lk]7ݮ���^�L�ɽ=�^�b��]������-��95�r`5X��4�!|���R�e:ʝ�
�u��r��F���@>�1���H@j�*as
����e��;R�+LY�L\�HxU��h��4��,X��9$gh��^�k�Ө �iI�}u�/�./��͇u>x\���*#�)&�\MwV�Ź��\���HR���ԉ��kASV�Z��0�����;Kfmυ�t�8x<�Џr�\�J���*���xvE! irс����>�]�9����԰��� ����x+D�&�����{�-C�h��x3Z{�2b������	5��,L��`���ߣ���ڲ}�n�ǖ�Kmh}"&ϐ��	țds�ݐ2���.P6�s[��ee< j*n+��M:�B���"�1���<�n\��m�ޑ�o�>5�l��ʐ��i��\���W�2b^!��;n�\C�f��&�	�74
����N� �Y��w Ƥj-�#j��~��kmɐ�,��)vtލ�;o��crA Cd'Ns,omb��w�B�����m�{�ƙj���bH㴽����,q�dV�U��j���}��Bydb�z�_�R6W�E�c��m�C�	*~��I��m�(b�ߩvw2ǹ�-�nDt�f��+;��DM5�^\&h|�8��ڡ��}�˾��t����t��3��Z����ek�m�-��픜�B���:`�kK�e�l�� �)��`��y�r0��Z���{j�
tS�nR���Sw��d��;jl_�s��S�2t&&Y�wӱS�����#����Sc�Kw{���38��/S�H����|fHM*��ݥi�R��KNjo��G����H�Q#�j��$-���e���E���C��ki���M<VV�5-���YI�iO��߹���,�	p��O�Ȳ��Ŕ��4�T���46�s'D'�`'@�@t��6h�Z&ڽ ��7��Z������j�H"�e8>3`�WGP��Jb��-`I.IxRn�*�7�z'�Ku�8|��P40�a�E��xh�.��VJ�&6}��}|��(���bFgӖ�l���4�����4g���ۘ՗߄�v��D��E�$:��Q�KV�\D��l��ĉ'j�B�����L�{����|���A�����8B�*��:д�P���)
��`���RG�������9�ă��T��L�M�lU�pP *�p3!:�����(�{*!��{��Dx�|���dHE=#$���?���'9��6�\o~���*F��ýթ��Nϯo�^�`{���2e��Nމ(�T��'�Ӽѷ�m�y�ms0�I��^B*��/@�л��,�\��a���hw2�M�T���ܾf��-�.r�� R�9�`�9����-k��}Rf�� �Q�?��8��V��c��}Gb~�!��
���Z�?v���q�M$�f���7}��a!_���+���aH�����i.\��ϒ�}�ڱ$U�p2�d�(�qu��U
��y{$a{� V�B�:|f�쿖ˉ��}8��K��M���u�;�����+ir�3�4�k�h�L����?�3<Ax�hzP�Ck/��[��O�7�q��!$� i1��bP�1|��)u���x��۾�S�ǜ����^2��3��"�Ӽ�`>�"<o��MX	
l��*U�.	�7c�*u�z��A B�@t��7�<h�Y��M����E�#�L>��VP�ގ���b�O���E���j)�y�J{������E��{�F��-9����ڮ��>�������������Q9X��=ݜ%����Ĵ�&���7����l����g����l$������3ޕ����~��ʱ��߭I4�s9aa4��E�� b$�&J��"
L��T�����ظ�Tã�[\����?0���3vC�I�98ڟH4Z=���'�cA�Р���S%�J`)k��Lr
j0}7Ʌ�'m̱����:���H��Nhƶ�������&��$M�e5cn��an�C��r��@$��b��>�8l�an�T�TWک��m)3N�Q����#ǥ�����ج�_$�$����9
H_Ը-__J�>�j��L�3����E����g�,�9nCh{���g�-��@�]9�i��+�ǽ�Ȧ��Bp���Dhb+���{�`b%I׼G�Cc�����'_IZ���W?��څ��7?7v�``$�kd�ވP�(��S&j;fO����6d�4ySc��GC�����"� ����}GiYa2S8ѴL:��@A���H@�
ZttZG[����ɹ�O��1i"��%���:YX�i*�m�x�?�n0'���j�<xmNH~�1
�\��v�Q� 5�i�����B�����u*s�:|0��?���e��
^�me�������]~"Y�j6�>���X%Z�8�M�R+v���TP����Mn�d�����G��-�6>N29�ĤШ���%���u/�&�ĸ�2H��Ԝ!&.n&��E.���O�W�$�;]��*X���E����f����a!h7U8L��g<
�L��M�F����������͍Lns�^�r�kل|S�J��P��Q�S�b3ic-�]r�-.ם�8K��OgN�p*'�Iv�	�2l� 跺e�!s�>St�ɓ�^܎h��������E>d��U_y�l�jɔ��-�`����}5�l6d�ٟi�d{��:q��&ʿ R�ąS��F�b���#j������N�����_J�89*wܑĸ��\�L��󒿮aw��1I���7�� �t�}�����#��y����#l�����2�؝�u���2a���,�lli�@�/�sb�c�-������;x�)'�S佧��L�{Q:Ỹ��H��ȋi��%�Ђ|G�k�6�Yۭh�j"#���31�5�/�g��ٴ�1�$�W���.�;��̈~��(�W�;x�fU�J��7mem�"N7B/��X�dh���'�1N�e��W��{$���|[q�y��_��~%�fu�
��+k>���z��7�9������{I�-R�o�e�0��j��^⿗(���#:i׭?��D��R�N~�8��+I$0)^#l�ۨ��`}:��#��ձ��G���lx8�y"G
f��r-N��!�Y6A����Pg��ʝR ���'�~5��[h�B���#$ъ����J9[�A,ױ�hz����4WzK�U"\�|	�?:8�=�Ш�/2ʃG�)oy���9Jq��&�w�������l� }�_@ܓ�@N�Q{�����4��?c�b��~�)�H�=_g�~�8���)�ތ���H��\��(:�����ϒ4ۅ?qc�D/_�?Ot4��6�[�k۪N��f����T���
^*E�%$������HA��㵨�,L%z'���ͬJ�nYA�i��,�ݦ�����Ҥ�#�ň�tII����v�D'�gX����9�j�p"�{�Q[��3)�o�{����X���*�Km��{��}� 
cB�.qI:H^�[J���GXb��7S7���e�8��>Mx� 1�&���Z��� EjA�2M�pa�n	|�֐$wѠ����>�`�Б	h��Q���^�`�_h��ב�����Տ�z�͘�n6"��b��7�Q�֡0�u��y7�+�6�����v��n���w�{W���$8�z��+J��WX=�Ǖ��RA3�`CA������C�Ř�?SqX{I�&&�r{���u����}\8��D�kX���\]�X�FF�zI�D�E-!��a?��r	�z3H�1��?)r�*���@-���"nD��뀼1y�Q���P겂�0���D�q,�VI5&]${�RX!���b�o9}����du���FD�Q�L�Z���u�3���� ����?g��^<�#I���A�Ibͩ?*	�a�
�Kr�.�Ҏ��o��Լ�]G�����+OU�1�)���do�	��}�� )ŧB��Ha;���&�H��q�]l�Գ�q���� XX��X�7WB���M�d&�M�~�o�8S�<Us�ȡ4q9���3%�Y���_��J�~�fx" �Ol���D�<�� К��k��u�vϏ+U��|�։N_7��U�0�5���5ڞ� I
�����&dN0���U��r�C��2�Iv.��"�e�*�$���Q%Eɮ�V���։(s��)���ٿ��b}��1+F3�]�F���5��ؕ��zs�i���m5��V���ç���������%=�i�9�e=T�UO���ڊx��6ܸ�fD$X���x���^�-�߿|�f�����<W6Hw�@����H#+�?3ӹhgv�Fu�Zg�O�� ��I�z/:�a�[N���\Q"Ea���o���)]P��R	����M9��U3y��2]8��� 4��h�!�݇>�u]r����f5��\!��w�3]��}?�)��ޜ��g�'��˶O�R�6�9�����g/�[*4zvA�Jݣb��g(lтx�V{ۃ��0y�U<���!�?H��{��abXJÅ�JQ���d�E�.�_���.�%Q��q{����8�V<!Xq�{��y$6F�w�X����*V�%�I��g��(M��\��2����w��E
)sC� �T"`+!�s�:d^����3��?���VE��&�`+ݭnb#�Y�v�Q�8Ji�w�~���HzX�:�϶��p%� 3�Q"��ߞ=��/�d�|z�uId������%�{�Pm��h��<�m��(��TQ���6�W�v�g���d]��Qs-��-;��6��_��u���ipc���'�V D����t�L��)�Y���O������I/��]��e푹��2w*q١��S�\�e٧�Q�cH��j�aψ�Y�Z]�02�G;�1�?F@9�~�b!mfY�C8"סg��Ή��ҝ�5�|����m���I�ӏ�C�;wq�I�t�
y�(����yb&�F�Ԗ]�����w�L�e����?�(��!#��ݩ���Ҍ|�)�����)��KI��H����X׵����,���Z��l�{�+~�����Axb7%�[Χ5?���Xw�x��h�vk�B��V(.��ij��Ϲ�z�jLm3v|�k`^&J�:ܲC�@����\v���҈���0��7��L��+�F���LU}lr��!��g�%��%z����1dr���\�+DG�[(w��V2�?���e��b-��ʤ�iG�-O��)�� e�ײ!�=۳쌾I�������7��3���2;��9Z����>ڐ�D)�mh��.zd3d	�Ӫ�N(R�Y�H�!���Ⱥ{{4
&B���5�-Y�g�~�Մ�i15A�|��Ѣ�����)$��]aF�$��|�D0B8�e�'4�X��5�䶟K��je$qC�a�����dl���4�a�ؗ��Kf"G����r>��x�#�뫠��J�:p�xZ�������j�1׉�p��w�%�)uz<¯㕰�5(�Z�UݽO�@\pY� i��>�g�'N�$Ղ���X��{�[@D�)�r�"���$`�e~�1&sA@0_�7��GGC^��2M(� j��U�}Bk}N�/�4��A�FC0�em2H�M��d�%����q�$'�����	�kv��C��|�X�ivc\4�aW���L{���M�������r>F���ëF�����U���f�_������(�.�����<_kȥSg��"FH����ȳ�|�Z�NJ�t�6d��JY�ɏI�tR�����CSj��/%-L����T�{��r���h�������```���&��Z�H��Iί3��
���xHy�Q��D��Z��_?^}}���a��&Z�̔��B�Z�E&W��>�y�ٖ��M皻���7`��p;��n�L��њZ����N�o c�T��N>���sTo�X����s��5�����M�oL�z�M�gkLf�����ԙ��5�ؒ~S��t��S*[�`Ο�� ���� ��I��V���,KK�P������%�P�O�6�?��;��1'�|f­�ц=y��s�[�Q-Q��86��K�AÑ�̘λh�_���zF����>���u�f}̘����!��X�Ξ��&�f��#r���&-Ł�0:���|�Tj>��ԋ���zz��9�Q��\�����������oF�f9Y������S%����?>���F[1����k�o+пpB+}���=Nt��:�%ϲ�WWݩ���!�-�u�3�v�m>�50�R
�,�I�y\�'�'пU��@b(��u�ɚ��h���w&�mY���m�ϦWl�΀{��n��	6�۲{�%�w�z�i_{b!OL�_H�>�Mpc%��s/�F���@��1����[�_j�0&�7N��%8R%����"��];힁W\�O������]E8��i3���fS���.�s����Bcm��2�\�tX|[wQ/���`N��� ��x6w�!����`DL�[R!��}�wXW�;Q�"�c���(��.���I�~���ٔ�\B���t�Վ[�W.T�g������,��9�����3$<\�������B�i�5���_�j*#7�d�S�ՑA���Ϲ�A�L���EG'�ʬZ׹����2�h����-;��L-����u��mϸp5��#56���)xZZw;�|�^��%T��0,4\1�x{Tc���4A��θ�m*��3��^���O�)؁ȠH����R��z�b[9�d{5��`_7��۩��.��񢧀`z�5�L��1��u�EF�Vg��I��k����Tes�t�k]sKLEFg^�Ņ��g�m6a{MD���'' i�]�����>���ƺ/a4{r�
(����ԭ@t]���'��M֝K�|j�5�N۝Aγ����Xq�BN��J=@�!��o��.�J�!˭/uW=�U�gM��41�B@.^���l�I#Jxӻ7ߥ~	����K5�˶�\�[b��X+��M�'�ڿ:����y�u���m���P�]l���У��6�Ex����ON���0jE9��B6P˦�4@Q�9W���2����X��7(�}r��M��B��]�T"d�b��E�-)�n��]%@�L��10��T��Xr�O9�apF�����5���B<`�Q+KO��/`�T� ��y!j��}#��r�f�B�H>�3]I���开JH��W*j��)BSb|���~M�fg�%�'t�*��ҿ�څf��W��:l�[Bh�_���kR�4��!��a7aU*ߍD�T��5��� v),,lf�sGiG���o] �!+O?$��o����Z[���q�|�dPB��5��Af�����VNUEK�7�9^>Sn|��a�n�x:�n��1x�oY��T5���ޕj�e"��*�͈��g�kb�o��eD%r�����4"N���`D<(��"��1��4(��]1�."�e���#�O���1r�*����þ����\��D�%�;�%O�|��+W��}�9�<�hx���ƌwπ{\ ������yTGbs�\�!��o5�/r�O�{\��Vɝ_~�����ZBW�ECM<-�pG=��\����N�p�w��$"��~U�mi�4�%�#�A>�����
Ue�o�\��@%��6�k�M�_zU�<�N�pL��>1�������a ������rװgxF�IߵV�_�,�s3�K&߳�7�p,A�u�y��ƺ���M'����z]�?|��@�(�����I�^���~��g�ʡ�fU�4&�^�n������)���"���G�1�lD�Te:T$�y�y.=E�V�O^���6#pAMq�JKr7�9r�QA�¥�Vʰ��vi�t��+�ois3���S� �=�$�xi����g�i4�o�L�\�j|�1��Ғ*��'b��$~R�`¼��6ȸ�:jw��d���_��vAWE:��FN0��~�1��	[�5��%HXqUU�H�O����\��Ҷ��<2m
=O(W䦓Ӎ&HyO֛O�e��~]@�"���H������Q��6�/���:W
5�!�s<w��W�@�H��ݛQ̓*�Ә��:�>�q���z���^=�����i��~�A�S�\$Ly��	Y&=�����#�D��?�Ό��Ox'�����4�u��.CK��((C?����}|��\�*�f�
��Q�9��Ɩ�7׫�CeY������s��<?��%^��&�l7���?��֬�)���X��k��pJ�AhPX�爔.�*�������o�G�m� $Px��ج����</V�I��'��yi3��Ƕ��줣Uv\'v�|_X�˸�̂E���G4
�X���8ɵ���D�j��{���<q3a� ��̍Ę��`�3
�͜�'Qɩ�������
h�Yē�󡕽l���k�~�(���8�=V~�m�h���P�	�<s��I�b� ��~cRvs�q���p�o���J�D�i3�i�a�@�.��[�T�ZdQc��)},�k� إr�HE���"N
�n�Ĭz��"���<+v���	:h��� &'G��y�]���Ģ�Eu���E������I������v�����<D�C�<��o $j��ї�Y�L�_�4�ߔ����֓�������4���[.b�fS�Qw�h%�-v7�r�ӯ�y
��>�Em��^��H�� ���gr|���7h]Yr�n��8vZ3���x���QҠr@�]�!�x&Cq�Ziڪ��� )�'��G�l��ن	��ߒ��\��)��ƃ]��?r�,���y�����l���1�zǢӈ�>��U�s)��;���f��e8\�ϿZ/b�6��9��πUID�Ң��J���'ϮK&U����͎4!N��y�:�BQ9el�:*�A�����=�M�<{*\:��� g?��������jl������(�Lߕ��*�����L��F�C�<n�J��3V/v��`�@<Y���%N[�4��N�GC��n�dF'Q����]�i��{�d8;�*05�3]���od�O�:�/��~%ٲR{�b`�]�Ed���!��`V;(Љ6{���
���|Au�I�F���^؁G*�L|�ۥ,�O��k@�[:��_�Z�ƛk̳h�ы�,�ԑAc�%�#��邠�R��A�~IAzNH�Rl��Ct��uNQo����^�$��c�Ϝ �IȈ�A�I��kj	ɊEe\��n5#� �v,���S!�^D�c�P�����N���M�Q&������Ӓ��������OG�,4a�Yi~K�3��<��j���Ҏ!cBmJ3t�¼Z*��-���@/1�����iAD/��F����D�̚��ˏE�����#W��K3�;�;����̻$i��ӡ��h�U�)r�:��Z�2��]�	�=��p���������]Y7AHm[H������@��;�f˶��}�7{ohN��s�܎�х6(���ũ�&r�ާ�R`8������{V�/�'����0�(�ޔ<�c�W�n�������t���G&�E��H*6π^H��i^ѥ����(�P;��<2�S�(0�m�9�<>�3A��*Qe4�����F�Y|I���P!f`����z\Ey���wv���-�Z�)�o��rT�3H�OG~��M��8��vU�dƻmJ��^���(���5J�@��<%&.3��cq�ƙy=[%���)���61��"��z`C���g)F��I�
�
{�HSwT�Ni�(�BsT1ND�?i�Lf�7Ð��6�'f�D����P����	,6q/9uoX� �~�5l����Y�"�L~R�����๎��NH�QJQ<i&���r�"-8��n���]"Z����
r����)E�	(�S������ϗr?p�*I1�Q��ڌ]A	)��5�c׍���u��������ZT#G�u�J��;[�r5���]t��6��)���z��9@���v� <㶠�/ �T��{�p}J�
����aG�GD1�E`�X�^Y�PW�1$�<�A����pY8��d!�Qg�F�o�������o��n���5!�/�M����#PH3�_��ß��;��׿N�:�i�~
a���fF�Gخ��=:�Csc�+�#m��? �d�qB��Vbh�<cR�Uk�I���4��^Χ#�#�(��(��S�[=8�1����i7M{��h,G��Y�LaB�zn�%t|�I捈?�r�r7ct	����t�����S|�:p� R:������.\��-j+i؂�co��I��@DV(��;��H��t��ms����D�����`��V��e��3UD$������0���~�D�ʖ[�+Lp��ֹʕ`r�U�|�R���R�:��y��1�`~X�P�
�<u%~#5o�kƣ���:̧�O0��S��Ʊ5�P�B��]h7 �$Mc?s���E�Y����a�Y���n�h�<���s�Z�ן���a�}�>���1b��[�����8et�g�?}2���e�DAT�ؖUf@ʆm���\��sſOLZ�q�C�|τ��C��3X�p�9�y|�S��ث~��,��(^����z�'չ�HН���ʹ~PB�^���1wW���Xh��(��7_�߁��\��>#�Le)�aJ��,TZ&���C�1ѕ���I@_�̣\p�"�y]���e7�.6HI=f���k��i�.�O)7h����#(9z�"��Ҙ� @dӛ��WO�|����m�qU�;Vê M��OLn��9昄��P�94�4�2�����6�ܱ~��Y�h��� ���c�Ee��>�"O�-_���|֖�	N#��pqv�MzPx��-aT��
u4�s�����.�C��t�'����h��#�*,��r�3W��mM���Re�`��!��osD��f�@<� �1��"+�.=�<s�w"D5e��(q鿍�o��Y�70R ԟM&�FDY���P��YG������ �8��h�.v���	+T)����T��	��W���-�W��{G��9�O���H�#��B-�� �j�Ԑ�M�ѴB�aD�.��u��r��Þ���c8�)�~��U.g����f<�����M�(۷s��ZvÝ	{~����N�@6��9K
Z�~�|���S��	�,��;�k�&��y��m�jlrP�P֯�Q'��8��>�"�K(#�)Mڑ`<��^���wX+����n�1wD������/��	��K7�¡����Ёj�(II����/`�2z��9dm��a�����.m�ѹ�
΀�H.n$N�k�*M����ޫ;�*o���PiU�;/��5���nZ�a�ա�jֹc�G�����zK܀���j_��L�3%�����FoLh�i�l |0�w� K��6���,�<�w���
0 ��#4/թ�xE�;E�P�b�LP۷�r#�dU��^���Ě<ѱg��K�_�{�ͣ%�Vw��:� k����P���@���0����ͷH
1Pm�T�e��3�֎�]�(G]�a��̹P�g5�3R�*,q�B�C���8���hF �J��F���8o�7�K:,�����Kx��r9ej���,PΨ4i���5) �Lsw�u����{~�9]����:�g�u	E�T��ݤa�Ϻ	������\ W�_���@S7�#�D'��e\}�8����������X'�R�.訳�U^.LX�����݈ǵs�&�Ev)�-7aV>7R֘ 8��0�QƗ�N�X�����-���[��q��0X���kk숫s�1+;%4w<K�[�O�P#v�zE�L`E3�(="'�XB5��ܲN]7p��N��5(r����w�r�	|O�G2	���ԥ<�0P5���2����N㠼�^�S�]?]��\1LWP�H��Ux����(�U kx�g����z���TH�6-�C7��`E48$����8!�����gpI�,G�ߴ�ڥ{�����E��W��a���g��]��0�f�\k������D��ޫ�X$�&C9�~q` &�5�"n�]���p����m���,z1�����u!���Ryr{�4�O�^�zMC��y6絨����2,��F� �U.�߬l�Z�/2��|���J��:M�f�+��:�fF�t#bZZq1���7�������m)�6q�*�R��m���4�hڠ������ˆ��G
J� �3���1�J�Q�f�l�L�.���o����6��S���r���ӯ���ϸ0��P�ܓH��M����Nd�l���=ݠ	��Y1�-�T#.�ay�j�n�U�#L�E�g�r����U���2NP��!J�?wd:y �d,�)q�B��kG��#��}vS�A� �^m�(h?�Z%M��b�<� e-�����*��n`�@���{�`�����d�(v7@���vm}����߬('F�k���+�SU�( ��;_���`�<��0	��L�M�L~��6���w����Sp��}Gt�_3�]���,�D��!��3�Z0$�?�� E0������4�+}��mX{y�����A�̒�֜����)�L��V��fC�~�Y��M�͠�m��iྮ��:Upl�(͘�p���e���E��Ȩ�Ʀ���`��0������9� �ɏ���!��r���7�6s"D��#��M �*�Wb�Fn����'P���Pj�A�&�M?¼�v1u�=�� ��ģ{U
��D@�ߓ5���ĺ"���,��	�A�/%��h�H"%��z%�v��j�1v��i�k��i+��UnK"����g�;����/�)<���xif]�xB�j�-��<���������~WHy��m����od�KA�
*jߚK���G��L��a��T�+7ļ:GBq�!YT���䬆�q�&7�)���'�#_�[�$y���
�.�9-�Q����`��!2d�x|�4��wt��k/`Ȁ�~h�i�Y�`6��S��B��k���d���
M��q��ld�k��=��"����|�f�r7T�qg���8g	�$)	��C��:ϕ^��/M�Z'���|������9����m���qb����j��ڙ�i(W���}Kpi�����r��I2K�ږ8X��q�iC�خ����'W���:����v�)V_���ނ��������2�ٶ0����f�H��zpn'"VeL��A�e�W]5�A��m��+aڠ�+���񴝩���M�R�9:רդ�f�Z����O��Y�yn�uq��Z9E����1��K�"Z|�)��yuk�D (ސCSM~n�j�7M�o�(��#��0��K��)��r{����8#v^����7�Ă��D�����`�)�)�{7i�=�&\/����b����.�;�OEC�ƻs�5֣pCӼ?�̎�7�?�3�KD���ЛL��\�+�+�oKI�fC�xeDU����ZK�@�P}���'L�o#�X���E��Ւ�����pw�jn��{눊41*p*�۷�܍<��3�i�/g�/�ъݞN���
\1����2��^>U���TJ@��M�u�����ߏ�-ϕ[�X:R�>%���R�A��/�R��������^T�%�nl���	��'T7!�휷�M@��(w4"�}��ϸ#��˜)Խ*����9!���MEҽ���q�=m��u��a�L
�)����=X�dȬ�ٟ���U$֟'@>R�(W�zP~���&mAe����g%k�I�ߴ�c�{�����dV�rmjI0-���^�4��PN��N�Q��]P��,�����tz��8�}I��!��,����n�:t�Q3Jn�k�
,�d6�D����bn�
IIX�����'�g�x0V�wێ�|)Cpk���츿a>�K��T�8�������e�=S4�Ƚc���\腆F�d��vc�JE��V>qN��qN�kp�+\e���0�I!jH��Ve�t��Z��Y�Kf�Q]��t�N���_�k1^�Ó����.��T�y=��%<f6���ʬ��ᔰ�4�磗�)��#]���~�"$F?�Fb����\�U�Q�b��7�-'�Iu��	-|2��0���ء�4V�\���$e��k��Z<�V�/Iǫ̘w�K4d�W�ȥN�����m�?�9&7��X�c� ������fSy�?o��2�����&�s�\n�'N0�4Po<Ea�`���Yc���Ĵ#�{->���9�]��cڟn*��sͷ���푵��aQ#�..@�H�ىNkTx�����Ճ7�ҙ��g.��,^%Њ>����w�F���>d�ac*��FA{|jy7�yq�xu@�t��ay8�B���iP�A/1�;�4�!�r��++!�~"�I���e�$Y�I�p7�z�A�bi)|��8Y0�״L��Maus�/1FĶY�=��nufr��ij�.���|{�5�h)�؏�9>[�/u�ٺ����L��W>=>��YN-P>}�Nݔ4�@�5^�鸂E����u��s@�刎�dV-�p"�GH�f�܂��W��q�d��%%~y�ZD��m��ls6"�DPy
���DiR������n��! D��wm�x�<������.� �m����8�#�^��@l������~�]ġ]���o�答���w��,�1b��G�E�-�B��S�K�Mн��B�P�j�VΙ_���吗�d�7"x�˰���	ĩ���hߏ?#*P�$�C��I��m�A���g8�R����O���w��8}���!mƛ��h�GQvO��*��!�����q4�����
��Ȧc��Q�GS�1w��*
XD�b�o��2q&�~{�=�aԽ��z�Vx��Whu�W��x�L��Cّ�[K��\��mU�	�>|�ٔ���K)�9M_ؐe
�#��؆���5�>�_�Y�.gȯ�/]7!R�lIv/���l7���G:S���,�M�-M۞:��y���1[Έ/�	�R)�Թ+=���\=S�>��Du��,xAv�]��qA�{���a��J����\���SÊ��>�.�)��<��w�0b�e/_�_@�$��9g����r% ��j�����k��h=�	ΫXOl3p;�^��@`��Z�ɳ�i����/K�&��ԘW�
���qy�.h2��o�<{}�_5���y*�>�S8�AE�!ȝ�G~��U �2��x�
�w��� ��|e��́��(�����U�Ҡ��$@m�NP^��f��B�Nŵ,A��'v5qɹM��&}W���j��l��T�G�Ee�I��~��{t������#A��s_���2��a�"�8bG6��������@���P���͵(^\�R���߫��bS���Ac�ޱiS8e^;y��60=�1*T�O� U��α�A�L���'�AT��s�����>mX�Jl���XRv݅�43"Z�O�:��^y�G�?L���$x?Ѳ����GJ��3���Q�*(o9!` � 31��)ş>����m���f��u?�T\������=��Z��׳��Ja8Q{s��rk�T������S-�o.��Ȫ�J��ȯ�@��:{��,;~�J1� �F�]$dں�yZ5�{py��Kbq1�]�Z�������n: �����5I�?�jB#�D�V�]�N_N�f�f��Mܫ����2��I��=�=�8�	��!gh'�#��@����ɑZ��أW��P�7���{Z�z�Ӄ�
�6o\���[)R�ϓ?g6�o�&�D6���t�2���[!D��RR��uм��ǰ�|O{�t��++_r�ӯ�Q�\�65����HFm���W�����RFc�,Qᦿ�.S��E�������1��y��;��r%�>�T���3&5��>�.�AH�Ǔ�>�����[/}�?PK�t8��4ԕ�q�@R��&��d���N�豴|ȅ��H�&9�b�1z2Xut���N��� 7i�b_�[ś��0����o��0�e�鰟sHW,=ި"�����<���xb���xh���\z[��"#r<���s%�֊�p�X(�yUŗuE�w�u�iZɬ�ۯ��g�kH�"��>��%ډ��"�=�/���r?��:��������Y��.��%�#,Bͻ�0���1�.�X�n셻yP2�7}�㐬.�>�;!{>~x���������{WZ>/�J(�3W��������4*�f>O>��u�j���~��4��`�ba�p+�r�a)��l��V�"\����b�d�]H�.��ݤ80��bSo;'Jȫ��O\a)�����t}+���.mb�2�3��۪3�����b���9��/���=fs,7�0�[A�@�oq�.��ܢ��^�e;�Q���رݩ�e6u�㋰�AK����������-�7�Q]p�,H�5�.�VuH�Ƌ�2�:ʁu)-f�&����}���wX��*�O�:a�al�C���۰�˸o�E�"��8��G�d&*X���<�lp��6��zZ8��5WU�|=��o�$�EO#iF��hˤ����/��*u�e���Ø��R	�(1�C	��av��=ߨ�Fp�IU���vIO�uBh��7��O�9���&����]c��J%��3�9�v�ڭ�(� B�0W�I�������(��<�u˜������������KK3��� ��S*���/=�9���Z�:��|j��=<j�y������ؾ�F��Po�o��P��AFx�['�O�]������Ge;Չ۹�lm��R"�GQޏ*����e�y��c���L-L2����>��Z	G��ʟ k�Yz�}�e@M\�zM�|7v����K���BI���O�\�{�X�]���C�*�V��	����}��==�}���Hx�.�$�t5���_6G)Z���W�Y��10D���_�c���jX�hD3{�Sx�$_Yw̪TQ$�b�;%�[C�u����L�=�t5*�j�E�Lv{�����p���c�� ��BC�/��ӭ��0�P<r$��f��-���1^-�:X�F��>)ɔ}�&��G�p)2�7n�84���^�+o��a�aQ�GL���o������c�\E��_*���/@��%���M��ϩ�� �;;M����8��q��f�������|�ֳ<��A!�&�R]�5xB���<�1s~H�	Y���q��A����:{�L���5*�����%/���ƛ�3�n8�B�`����-�b��`�Vr6a<I�e��|w��"��|t�	�1⻏Vت`��z���O{t��Ի~u䭳26cߠƋz��Q��Փ�4��W^�97��%O�P.*Fbv~��Q�8��P�Ѕ^�� �E�B$t�� �+��F��n�2 �Ɓ�{�M5J����O�E�ͭ�
�[�Y̐i3��H�G�7��![
ϧK�N���3�E�f��!c|IT>��xbq��}���N��<��_m������-�`��#3�����3Z��-��Ndw�`��g�!H��;�9����A�����80b��*�5)<���b�K����� |L����/KF$�.`ڀ@��D�V�T�#�p���i�l[��'a��W��N��-P�p�жjҖ�X����-�3	���!�@�i�_��B6[+>���H�S�d�(�u�5	�҇�[[������Cj!;ax��aZ*Sm�4	l9��r�D{�FVfݗ�6�;���x��L� N��A6MQ���
�ؗWu<�"e�h��Վ�Y��p������R�XT��M�6�p�u�l�O�L��w�=Yh�v���N�T��G�t����5�  P����T~��>�A�R��"�*n�Y�e�&��� ~�6H��(�����?�A�͢&���v'q�-��,�f$�q�Xf[��	�Q`xၹt������?����Jӣk��8��a�?�C�Sd''i7�1���`$������5�Gbt�w[�n32`gǗ��OѲv�H���E������@u3�r6O��R =0���%��>*�J=�j#�ٻ@�&��weVvibԐ�ӢL���9�]A]<E[=���.M.�5�?i��^-P��~J�:�l_vE^G��˟2�kT$]���n� Ӱ»�}�ý��]�f�f���x[�37Z�@n�օ+F�)S�dԔ)#�ԅj��N��"���s���"��Vm>���>�L���O"��'.:��w�vn=P�!��F����ȱ����.B8Pr���������K_�ok0���`�O7���D�co/�b];�����%):eoUҠzhDZ�a�	^L-"�5��V_q����?�q*ol�j�=��	�n:3b��ȥ�lDZ��j[�­B�8�(x������_(G��#gjDu0��Q�y�E��hˬ�����\�����÷��$H����K�J��B��F�B#��F���E<�{��(�\�n:)^$�VjV}g!�����G��^�fK�EB�tEfTOǅs9/Nf0	�����ڀ��,���ϴ��(ӞS�+KK1c�8��g���!Qf}^��r	������Y���r�`��<�ނ"��Z1~�d���A���?P�<۟E��a�50��"�N� W�����V�&MWY�`�!9���}��L	?�j<�C̥�D}U?/�&��n��L1��h�|�4�&�G��'�Jc`%ǵ�Ν�(f�r�6"�����y钠l��b�;y,>/��8k���;������G�~��k����n0�Ê����̍Lb�9��ֽ��m�ͦ������6���4�!ܛ�����xy�p4�j� �����e�9h1F~�����	�%q�VgLb(D-8�����ϲ��g�������g�ȑ�������%9E ����8�q���/�_����).#hx�DUn�1�(�/�_�_>��ٍ����1ۋ)2Ur��*ځT.kd�B��ّ�B5h͔3LՆѭ+��Jje΄��/a~Z�9̿��ƪc�������{�2,�0���0$��ԏ}�~���Z������h����A�|`;��3!ɼ
���!"��k��	#'B��W��9�SG���w���mgԫ.�}]e�9Q f�(bw�.J`�n��7�_3�S9OL�80�h5���?@C��P����e�C-�״ ƋzL��q�1c�u��;�I�2�{�I*�Қ�9"��ћ�6�t8�^�
��@�w��m�V�P�Y���S1��(����.�W�_�W�Y��|����,8$R��F�-�l5���+	t�5s�ߝI�>%r��lJ�� WmI��3k����������l�J2Q��;��y�V8��LDb:�P睃���W�*��f{]���{nA��4��� ��vh��f�[}�$y3���o�Z�o�|�"�ІU���������	�I��7�*8h�p�ϑ�n��r�B�+�����7�X��dSAρ�C��$ȩ�C�Wly�V5Q�NRZj`���(�7�~:��{D/��l)�Q[K������1�:����i�����ڵ�{0Q� �R��	)U+�zX���R�I�#��v�5�{X
$x8�c�[�ߣ��z��'2}&s#�d����j@�T�7z�=^uj>�Q�Q���ak�i��fcd�Z�>�Fa��B�,O��V�[t�Tn6`�_���0����nx[1���u�j9TM9i�Cx����!S.�n�ݮf� v?��������w�)_ QWX�0�N��k�L �!�ei}����hq!O�����F��̂ ����ӳ�;���ʬ
M�҄��wR�T�\j�H�C���V��bz�Ċ}D��(��r���[@B�U�{z~���d�B��eJA]Vp�;W1$H��PI[�}^7zS�6�"��6���;<:j�有�Uo0N���rh�Q�q��y�+�o��{F�{�����ǔ�[�7�ߋH
ݚ[r�`�g��@�.��0[5��P��@;h�ǻH_����R�ȵY��Mط��FV�G��˃��;��KδY�v�a�Wڼ�� F�6��Ef�iH��(>l��/bC��&��u*�&󵚫ӑ�j�>W��kLX�t���$���d�A�G�5��πD�?�h�&�.+��N�)�����$�]�	��)�q�ǉİ�}DK���_�^.���f�c^kHY���ӹ�.v@ߖAS�� ����WƯ����\�Cn�pI�W�&J�G+�����@J}���k*ȑ,W�ذ�R�V�&2:�3<�2��߱h�~Q��l*�lr³�پ2:�旍8���5�Ѐ��[�D
�[����W�aDwX��2R�����;�2�C�+���ۤE^}�����r�x#��8��V5QJRC�Y�|bFȴ?��	AH��}� �ebl[0�B�f	]{gt�d��n��V�@d���r|��*m.�l��`�eC�`�Z�W��=���"�3l�x���Dbێ�0*C����,sk�g��GL�e_4��<Iٕ��˽zұ�qï�pi��xɣW	VM�R�0<���O�y�Q����l��\:�!�q���У�K.�;�[9?�w�$��ѭ��WÈ4r��At@�c�~k������A�K�%�k�B�T
�wnڪ5w9�A�x@+���4�?�W�N�S�(�ݰ�֖�].#c/z3?	�-�YXV���{;	>��Jgf��O>�TT��8UT	��_d�;L&�T��@溈�A�Y�ڄ԰���6��s(��Op��$�횯E&[�X��n�-j �bG{I��|+��l���7Q$O�J��}f�k����;FXȡ�7�aY�K#�k�V��!�f��6�SC�Ws%fdH���6I1z����	pS���� �n}���c$Ec�'w���nS@؆����K�ތR�۰�hɍ�+�\�����.��3�D2�S�\��"C���ƹE��5�g&���F���������&[�~(i E�YS~o��V�'�(���ۨ�D$=���1��g��M���4.���ii7Ę�}�%����ˉ;��Ы$L/����"(�R<W�0/o�a�I����̕���>�f���C�wEm,;��`��D�������B?S˥�Lt7��+��h�����"�@��v�����U���w���,d"/�FA��曽t6C�י���2�B�c��5q�W@�)�pt|��������3�Ҋ�~�/���=�<�N�&{y����6O�������br�?�~)��lL
녠��ɇvo��~�;ηa(E�{d��Q.�fU��~EX��!�����}��`��$�`7�|�c����<���һHT�)��M�3똌[���L �|�`0P*��nn����j�Nug{����ل�x_cp�6z��;vWd�Ɛ)���VTu�09x�Z��(Jo^�o��aM����~RZ�{9�rA��I���{�UNG=������̴墱f�n	*���2Y�p2���@�V�5Y>�Jv���s�:�>)0L���]c���i��*lj="	��݄M].��>"���r'VM�:*q��괩��ϻ��ԺLq�t�+#Ư��zޟ��4��^�L�H;-��oΫN������Z�6fO�gcf��ډT�ܝU���"���H�r�]/Ӊ	�q�9s{A�w�07(�W����̫�1���W����C H�O��������ơ����J#FT;����Ʃ���]�/\�c H`�K�r����F��8AD���|n��@s:�Kb���Q���T�Yz�]�+?��?�Tڨ���G�G�P@:*�	A�0���r��6_84�|�4?�df�DPڤP�A��`�+�{�9C�K�O��5���n�[��j����)������T&E�2�eZwa�ΰ�
M��}�����th'T^�?�K1��b�őf�a�G�dZVf9�>�r��M�᝜�h¸bx;��NA=U��
�3�+�qV-G�g�	5PQ�Sti��W,�c'r��'{�����^���`pA�<���������P���]Z� �?����5N�$\L$y���˓���u�j����M;U���͵E��v��0�A��5�E`�v����F�9�2%�0��	�p�ƫa�B�)��rZ�_v�Ƣ�Hb)���i{##_ZF`X4����6�8̎�6I�$�>^�>�	�Ê�����U��7�e-���	]��t%<\�E�O�'T
i�J�b¬��
�����'/�C�:	�HŎ�N����籚�U����`L�d��h�'��c��L�l��ͤÙ6��`�p��3��b�qF%[��naY3>�����q���>�w��/AYf�@��� ��|E��1��~����N�sP��q99��<^���(^�������x���/����=X�Nؕ��+,�6*浴�͓�c?�b������d�a��s>�~��"X�@Q�R"uww�j-d�?�D0H9_���۽�+�9̊�i�a>�aٰz�������ֻ�2ͧp>#�+*F4P_Z]b\�ކ� FO���<�_L$���
��˝����h�#o:�W��P>:r�o<Z�4��	��Y�kg�n�o�}R��s���)|���:��-���O����I���#z�  v�7@�h:�r4/��)�$����nĿDih����	�$���tzV���S+:�m�ǡ�n�*��\Q�U� �R!�>v����Gj?���� �;[��^����ff��Eh�%F`ֳ0Ig���%��w����c�����Ô>5(��6�G�8}�Á �	W�s(a��^FN�K�5�! � 6ϣY��<N�K5-�%x��b�ôN�d����O|��bX<�+�BdlE��S�37m]X `�Ź�6�2"v��]����*�s@�7O<!%�Ԁ�3E�nm̭�� -{T�F�������>��Q"���$>y3�^Zf�:�k�V��Os�A0MkU 6S�G��_��	���?���J��t��6C��6��R�W�-�q����d��	�mM�7���D���v�#��� D�2N��Ľ���[��$��Wʎ���Z��%�8q��1T���.�X�8+ܾ�Q���S����z�/�%��^��Wkై榑X��>@]�9iu�]���lk���L���f�2��%�7��#�?��	ҎX��K�C�
\���Nh�.汐���_\�H���62��z�4y`<�������R�y@2^��R�TU;�Jt�h�26|�[���+�d�kL�vL��=�}�H�ُ_Z ;E�g5Ϭ�iIl[�Z?Y�Mn�v�߸̝h��fSo�c,���,gD��NRE����U��Rf�
�u%�E�]��ɍP����|3��3��/�D˹8��D¯�.SDQ?j$^<�גU[�i�J�/<�>&�>�'��R�	�:̣Y�
"�����7D�6��I�?��ʜ�x�!��A�l��
���?�h�ђ�~9<.+� {P<R���t ��UM97�A(�
Aպ}8�J	��a_>��H���s�:�f6���-��"���;���<���A�s�/��g��0�.���%�������;���\��]�`Y�8I>�Q]���1���bZ�_ǈ���5<䠙)���nkY�k�(ǻ�t|F;�Ph�a� ������i'��bI aU�Ъ�/	��,V����~�|��ۘ�t����^�����>��9ل\̡#�{�/���옱�3E�Y�����_�1��	x~��ҙXG����n��.@3��|<��yl����cX����du�&@�?+_�3�z��<�6�!��'Y�ޞ�9��G�����W�U�^�����J|�e��I��>O9TK�jnfZ�of��*�ⵄcZ���6�]
{����A���Y4�g��o!>�z��Z�p�
L����;�K༻D����J�7`Ǧt���j�93j&< #-	셂MA��=͜������n���6#H��n+*���΃kH�#�f8$حY�	���H���ڎ?OՍ�W�>^�:���ra�ea������T����V1�Ut�MB�Y�N��#�߳�me�d���3��>�rXY�`�Q2���I�������p��&PG�'�1�ubQ'�kL�i�\x�,�z�T�R,I�vA����2m�����Q_ֆ\r���L�V}�@��� �-sg��Ьb��HA�&,���sgǂ�����3�X���M�KT���)D��;n���lq����5\؅Ww��?_��VMh�������ZPX����D��o=}�tP�x ����斏M�D�qzA��Hn���Sd�.d@�j�/w�w�rm�g3���t�e��"4�ߋT���gz����`���Z3���$k��&��� k[�r��i���ׄ�>���4c��#i���3���(E�"����@X�"�E�d��X���_):Dgay������X���c��^��t��s����Y��ԕY	�x���ӱ`��*H��v�#
]�g캯������*!�o�<�J���9q�\f����ה�汅�Y[ى!�%w��Uj�/r���7�P�u��81�#��k'�j�������V#�����M��w�8#�t�����3gYV0��{d%��a�%@�76����>�>2�ܷ���DdE��%ve�~�)�����Z<bvD�]L��묓L�zK�t@��4�RH�$��8�9�`o�T�U�:����I��|�],??Y��Zl��}'kV��¥Av:��=�XF[����}�U�g���mǦl���K�hC�kN/��ce7�;���:�J���?TR:�6�C�@��d^�y!C���<���z�%�l�7hb��G*Ѓ/I���]�n1��mg|uױ���l�@�>L~��&2 U����(��oyV�u���kQ=Td
����X�q
��d6��]):녷OpG��_3�z��D����ˆ�O
�����Fgbw��u�\�2��pGK�V��t������J�1`�Cє@]"�f�����l�tNt@)H;���L��������U�6��_
��ƴo=��F��J?w｣$�I�F`f�%@'D
L#*Ƭ-��vB���B�#���E�~sP�ڝ����r���T�
��rc�j���_��垵�3��i6�]�k�ђ��f���{e���xt��z�c�	��y�{�T�tϾzK�������7��0��r�E��O�X���Q]���þɃp%�Pai�]Q'��V`��<���ސ�
/$����cĔ��|}��V8��%���[���
���ċ/�ٙH}ve�G�9p� FVu����"���',�"H	G
���k������8@�zr�+��*��c���%FhK��,�!p��ˏFI�&g����Z��)Rɧ2�5���I͸�+��z_�tx�V��_�2�)e	X,�����u���ĐSpq��1��}��
>�iT��e�C4�nz�Њ�x�|fLA�{#f�]M���m��׹5�Cr垐DL;g��)� ����_��INw���5��Ҟ�/j���6c<dᅮ)����&G�9���	��.]Y?�r����3����Gb�X��։�	b��X��9�I��̘��%D��s���!�3������>K'�U)�>�꿍'0]�8(g��]ʎyM���ʈ�x/������>	AB�����^��}R0�Ȇ�43Eh�X�z�<-�e�f��}Q��4Ĕ "�í��}ٹŜ��D/ qӆ"�5�a"z�
=ʷF�qIH"H�̘�u��Jֶ���feM����2��GHnưs��j,J7:G�h-	�g�h�i��3�n���P ����A;a�Ry~�����ǹ�[) ��1�����keH�+j\�7(��ݙҘ��
ҺawG-`��|*Lj�Q�oa��Y�C��9>Z�Yu���*E_b@Rב��r�읍�3�a��$��׎�64IK�܌^����ghX�AW�]��  :�s�iQ�60[aމ�T���T�	1����ɓ���1U���\�#��R����f�Z��N�E~�|�h�S~�4O�6�HYE4
=�Gן�4���Fqٿf���K�V�0��>|�������n�f7Z$�n֐�@S�؜W��iIy\�SS�P5�w��d���E?�c
�LYD�Sm�8��H�fbħ�)��)\z&�4gc��BU� ˥��ӳKU_�
F�D��-wt�����XX6ǜ*�y$�Ć��o��d�c�.�k��s�?
��B�x�^6�u��Ip�N3F>hTß��r"'��������R�D.]��tDoh�~���]�EB�&\q݋.p����u��� ML�|Ak�dd3i�s�oi�K<�K 0���ݍ��Ԉ��u����G?�x�����(�e2ۭk��C�Z���`�R&0��&�y.��]��Es;cI[�ݜ��󚴽�a't���x�<���&b�w��:��2���8%�܏�8�b�A䌛��9���0BB���B$fM�����1�G5]�)By�����rQ���t�����&hZ��?��Z��+�J0���!,��V��`N�k�؟ڱ�k|cS.�b^F@�/彝I�����$I�aW��l�S���t����Wv4m�G|k��'TEɢ�5�q&:>�V^�D,O+&%7aOs��g֑�h�D��_�;xb=ė!�����rK��Yם�۵����]�sS��s0��+�;�������8;�'��ڛ�%�F0��Fp�U]pi~�qr	tX��������+ks��Թ6�6:b�6����N�1fAW����P킱�����2C{B6�'����F&�ÚM��h���;� �+)㢯��Fy��F�F�մUC���>�i��LiW�����&�_��l���.�����w��/"{Vr�:)0Η�S5����Q ��9:EA���d|�15��iP%��X�[F�B�R^c�/�����|s�Aq�>�iQ��g-��$8����oɠ���k�i/_3�2+ u�`�^��'!�\
7{���5����Z�i�����?h�����c�^c{�>:A����9�x�:�X/BZ_6�b:H3�!,��ҷ3��t�ɿ�m�$h� ��cn �ӹ�J�k\�O2^�\d�|��E�X��"u=6ϗ ���46$w�Ȯ�n��{����kq_�KYp!Jne΀%����=���%t�$������5s[ķ>��H��G�V6 8Q��,@PC�Z����Y)���0E�7��F��o�<�($�<��Aȷ"��y�O��Xef����^$P�\�F�:���f[���1�����ȔqIW�R�"SRH��0��3��Ci��K���0��|�/��s8��S꽨8TN���Ap*+��]�SEM*~����k"L�KqX��.��fCo��F9ŨP�~�K^ȶT�"h,0G8='�� ��aF�͎n ��,[OARC�(�:��Q��-�9W�r� ��#�hzw,5��u:oc^�$ŝ;���3Ɗ%�Z<�S���k3����U�k��*i�L�G=��	��-|�����6�9�r�gJ+vE�t!�H��.qn�#<�H�'[��F<\6�{�Z��K����q��J�0Tl|�oPq�B�j�fн[!�ޜ�
�W��'��1/�6�pb$�>�W,Us,k�.5� �)�d���l�h��
����Y;�f�)�-J
A=�5;l��PQ���"�#H<�"���;58a:a���o~p��i��1]����i�*�O@F����M2_k�|"'�Z��4ԬV���U<dC��F��������5!�E��=�0!߳=��ok �E(V��_��ȇrK�Kc�}&�9����T"o��hDh����7��D*I�:��$s��<c��+0LQ����ɲS6t�ݸe�`���a�~g��jr�Oa ,����{�x�~e���k��&N�g	_BS���Ơ��B�#��7��ەo?�D8�ɵkyRu�i���ء�b���!Gj�Bs���a�N�\�]t��eiOG�H�R��c4�%~	�����#{ ����zBr����ITR���(5P�S�@�V�o^�?������NkV���3�����Bf��R|�~F����o1�%Q�TC��`E��ǻιl��*ہqŲ
 �_�9C=1�u`���L6�XǶ��3�W�"�����=�<�34S���@�/K��lX��s P�l]�_2fo=��i<��d�XtW)�zeP��x�e��O��g��T$Ky�r�U�
��(p'����!��(őv�W�����c����X�Pe�p槵k5ZA2ٮc-�	b?�	;�.���A����h[n
��ƾ|f�E�`��N3L�No�5k�Tg7�1[$�ZA�e�'���;/i�ܱ�UpW�7ݎ����v4j��>�3�w!$tqe6��S�䉞��W���W�Z�9�:�V�8��DrUF�H�|��^cOD�"��-Tf�:�y����"'� @�1"�9��� D
��s�8F!s)y
T�s�&�-�7�����K��@d[a���Y�&8Ȥ��ȁ�r/���m~������<5	&��XC�̢�dծe<��;���Y�Mȱƪ\n��dh� l����cş�����/>���T���=6�s�'l]n�8K*�A�上�3D��.�k�p����~V�98��&`�z���VN��2m����n� ��[��o7<�xU�C�J�����Z�$�W���FM��8Cyy�4�E��#%�-^e�T���|��x��C)�s$FCQ�b����,����h�ڹ��a�i�M��$*�}v���	���r�!`9��@⥵ڡ ���  �h�:�w�MN�A��1E�M��D�1<�$��p{��Y6[l#��	�u�P�q��,�=�E\����@[�kO�jt�Gz��!߭��Tm��a��a^N&�5P|�[Q�4�	��BqM,���@����U����`���۽w��i��T�H�zͯ���}��b�';\�0�#� !r��'A��$Ր��=X ���U��>q]�&��T�Qg)�-���*B��Ҥ�J|�18�CIf] 1�:��ҝU]3ӸL��|���3?��#�@��A���$�;"���p�(Ke�sKx�!���IZK+�MvS�{�]�J���J!���-���Q~��3����&�����,�H���c2W���p_�0�x�5�sK�Ԋl����iŝ<�#j݀�\�姲j���g0;w�gzz{�le]����(�|���4���%BF�4�VuÃ����4�����]�`�o��rDv&"���%C'�R�N|����9H2+���>�ϳ���<R.�P���Q�sG�=q0#�ּQ]��Z�*Kk��G�.�y�MGCYw?�n�����R�ߢ�S������?~S|��wsī�3&����\4 ���S*�@v��'@��*���]~A�i��B�,����H4z��zé���/��	�Ϩ���ʡ9��*��(��m��k�G�b���p$��T���ϵx_��Yq�l+���΃��J�/�U�{��H�r�G��n��Z}�Nh��Z;j�ǳ����W�"E/X��ʝ7Y��+\�y�G� d+��f?��B`&(�N�|���пPr�����Z�0�|��pj�2��_OLl��E��V��6�w��t�vR�Ic��h�[�'d�cݦX��l�KK��w��lck�B�/�A�5�&Ty"��R~�_� ���� ]�`��}5hU�|&���������X���#�f�8Z)4&��\'a_�@����"e+Wö�
���J�kQz`��1Q�ҵ�r�M��>��xuPu^��Y�R��ǟ=�{/ƹњ���-��f]~;
~6���cY8�'��U��T��#��uYn��`�M�~��q2��C��svU�����Ձ�=�K�(�Fdk]���)wą-���:�Þ�E@������s{d� ��e��T�{r4��:��֕S�Z=�S����ɗ���
p�����_4`������%zy���m���+	% �Ō�;48s˯��i�]'�20�V���݁gm�K>���O��	T�e��{nЃ����2��"�7�B��ތ����[�9&�5�	T���[8�G�S�$��:��ބ.��}�<�X%�%�P&����6���C�o,�����˅��M<���/^^����>c{�:s;`7�~������.Z�S��	��NC>����nb������n-ָ��!�&̙0����]��Nf�賟�w��j/RI���(�衭@PQ���t��G���%q�5֖k0�������Α��/x��1�ve��lE���7��걨vň��> �¿��d�U�)�e@��ថ���y����A�(d3r��lY�`��&�$�����o�ɭ��Y��-����J�-������l��KY�$P�uk�'J�j�p�H�d��#�dF"J�~�%����k�\XV�����t��^�Х�eEݰ6Ff��V?�&}�j=7�}k�c�V�ҟ�_;n{��a�*~���:�?��<@� ��w�-P� 4�7�fxsi]{`��Ed�<�w\?I�/�ÕgYw��Ѫ���o"�۞V��/ �R��e;P�P)0[��0$S"��;.�8z���F�ص@�GF��6jh��h
jKc� -t�W.x����ܡ�	��nWj;�՚�v����^��L)�7���2�����k�z��L����h�k��֚�O�}���:ҁ��JjҊH�!P���g�c��տ9�7��5൰�8X$�o��w��h4\��9�To����䡈��G�M�K-��3�o!�y����d���*� YL�mBCM7$&��@R�ò���!z��zXq9
O�Kv��Ϯ.�תX�AK�*C4��M��k�D�K�#
ޔZe�O5�H��ʊFm! Q2:�%ʕr�Vܨ����۔�"�~�tg��ڃ*����	ܪ���Tݣά� ~Cb��#�b�t�OdW�A���X���1��P��4�B��j~pB�N�y�s�?ҽ����J�ל$�t��7�����aԨU���-���{I�Ji�@�0za��I|��� �Ul������U�[v/�n]�Y}�R�Z)l�, �@�2ۇ>����IrM�����滁��	 u�@�˗-2X����ߎ@���xZ���%���g�����^����� ��ԁ���3t��U�ؕ�Pz����; 46CI}g��ԕ$�ǳ'\�"���-�8r�<�Q	n�b@�����Y~>	L���o�r��F+�U�?~��g�[��-�	Xn���k�L -�QA�Z�p�P�[s6Z���j�&e<�e�����YO��\{�q|���0��lAJ��̈́�3��TݦYzx�FJ����f�!ψ�A�~��{�?�[����[�/�X���֑+6Q�h��Z�t�I���]��|.К�+]�����j�	��[١g&i�����1���e}+k4xҧ�����X��2ӕ���2����XG����S��K��7�
�(��7��@ȁ�5�Xc�����:p��{���铃d{�y]��/Y�<P]θ����-����,hG�s}M�|��%�R�+ۄ�����&�q�<Φۀ,��Q26��3� m�w4�Ω����]�)ΰ�Z\�b�S~��.���^b'��j�iԁ߿P:��{��D��.��'�; ,��'�Ԩ1p�^�n+��a����߂R����7B�[�J9*���2g+��h��Y���_�>T��I��J�J�����r�l�T���j���x�E���-y����H��k�&�Uy�Ak8��������q���ȸ��s7�<���CIPciD�#�۞�!׋*G1f��v?8���*q���-s��Oh�F�W��p� �WQ�`nv^�$�)��\�ޮ
y<z�u,&����娲����8�WZ�7ڎ����R�p	:�b�ė�N)x1���P-T�O�5�������׽��xg�V��V��j�[!���A����5ZB��L #��v$�C�j��B1�����u�1��-��A�������=�
Lu���4R-���6���W�hW��鴸�|��g9LFq�(�,�W��Q���/�b��w%+C�@X6l�*Ʀ�z껲�΁��iH�@h�4Q��s6;xǄ�-GY᪞�uy�eK��7+����J��y�d���w�e��M���!�?���=��k� �Y�%��L���'�8uw�W$��ȯ�qb^AZ�}J��������C#�D������߂��9���U��A^#��Im	��$�K�Dj�+C�a�=Veޒ��Q��w�t����kZpIb):�t8w��Q�4�D�@$���ʙ��6V��sMݢ���i��K�0Ax���Tى5����Mkw�&@$D�VE�Ԫ7Q�v���#�E���0bI9� c�R%X�p��B}�/h�F��O��moBO-�āe���>�5�t�JlX!I-��k}3t�9�at�W��vg@!\�&����ģ�K���VhMEJ�	�b¿�3���u%2�8wlK��uQ�p;�Ƶ�͸Cb���;�+�o�\����TiK�6Ip���	���y�^YFE��fRx2@��0�)��s/����:�y�Dً���,�܄/n��t�ܢ�ط�u?&2��jg�*y%�ENtu�����AE���k�@OX�`��?^�GA��_o����XL��M�C1j�����o	Dt�!��M�1�X,![��d-�ţA��9�����1���L ��=1�s=�@_�y����37��h�'�8�/7�x��E��C��KAyl����i��j���ՅZX���z[z�ذ�������i��F�؄�9ս��|~�e��G�OQ[*t�a)��<�����__�,��nq���nR)�ш	����Rg�W�e�ײ��PK�~$f��)4��� Ω����I̒q�W��b�p�.D�G(��I�@<���+pJ2��KQ�A�_����-���Q������ۙ��<ن��]��O����P@3�rV/)
�\G��U�6�[�����0�	�L��.����<��[O�����A>?���?�G��ӓm
����k\�V�cJ��y�N�&�A��VE%���޸�=T1v��3i�1��A��7ɖI���	��IYJK��hb�d/�_���#k|�:/���8H�W���jӑ�vD1C2uhT��B��弛��xG�x4NU�F��b4i�
y�m�ԋ/��B{`�d%2Ut'Yy��zv9�d���Q���%]�b!��@�*T� L�g��k���u�G��c�Ѯ@���^4n�G�$OaM'y"�y�Nw�+6�F`/���e�F�$j�ë��DtY�ɕ+._��?������L�e�O��,�n�U��p��CqW�)�D�]�O����?��/�n�p}s;�A��=�<)���K��;�s�5S\�'?��'��a�Xyאߌ�xg�Tè�J%O��#��.~��H��=\4
���?�N/H�������ֿ�\�_ o��q���S�8 ��B�	��q���̘F� �sd�QY�`7��%����W#&����������QkZ�����q��k����d�]����W��ȧ�a/�m�'f����P�Iŕ�D*��y�?����f�%�����^�"r�$m�a�m���j8�	�{k�J"1�^�W̑�����-Wt.�X��9y�Ԅx���F2�aF�ݾ�;,��n	*Ķ(N�_)�Y��J��_��,_S�a� �du�>hq9��rCh��`�aS����0]7�,ݞ�G��m[g�j@g�q��̸�8��k#�n �eZv�cAKe6��0��,�H�szkhq�Vvk�gg�S���0M��F|+n���+��^ge@g�%8����.������0Zj�G�ii���EQ��ar&��b[pA��~}�>!��v�v1��:E����n��<�#�B ��+7" �V����`��w[�=Y�I5v�¥d7���!Lk�{&!D:��9dE3�O�S�����Βl�俒bڄ�l~��#�
�kt�0��b�4�����`�LR��Zo�z�m��_ע
d��Р�"ރ���k�F���xh}Z���guW�a��g��+�>�58�쒒������7��U�s�$�έ�ṋ�]�U;�<���_ܑ�Cw��ϯ�/������J�oF��Q���²��7�X�H�Ӗ�IXn�8�&�����oX�B��L��4�J}H��5�˼�զ����[^[��7����re��66���^����8L��c�N�dl�iG����B��g�C�~��t��:8��A��A���\W+�4^%+�ji�N��gS'M!�3�Tq>4���tg�~�^+�[�?��@:Au՝WT����0�z��ÙS�*����ZO`���<�L�T8) �'�i��~���O݀�s���̕nA��F��_FL\v���e�g� �59/�5SC�W���d"���862������e�n�Y^>�.c�,d�w �Y�\������ ��yH'����]1����d@ x��8��[���Ë�Ew2��R�G�`��[BPyX�S���y˞�U��|�w6���zk�H8pOJΏٝ�`!�4�29¢'��\������qRF=g��0�)�0���2|��3ݓZj&Q���u<�3[zL�G�wـ�n���S:!H�15@WK�����C?�[�ܳj��y��eǙ�0f�ɏ��'V͔3	�S�5��:��@�~��"[��?	���`>��Ҟ�-,�%���ǒ�ؠ!|1�a�̷.'<�U��	���h�:��wIA�FWU�B�]Ȓ�{_�=ֆ�%�-lY�P7*\3���g=v������m1F�=���0�֊�e? ������$��]^jpr����!|��mB-�`r$�Sd�S\ؽ�@b	6��	�ū�N� �0�Q��S`�Q�8Z�ӥ��Ht�u T^~�"T��Y�־�3"����/-r\�٬��2��G�߆�7�f_�Bg���q�wR����-������6����h�vD�����:G�z����m��@���o-yXcw�x}.#��i�N]��l�-���t�Gc���5:ݶ��ZA�'І0��F�����zH��٤��Aᎏ�{�KW��_��	���$:w�k�����bH/�U��3�1?%��G����:#D�_����1%��c�ӈ��-S]��
�(�?"Ż!����>�,���A��.�
�����GA���qR�N^�hN��U`����$����uh.CW{�0���AԹB>���L�_e�zҊ�g7:bn��=>:_�I �Et �5���â�t�����'H���Cu�]�����w�����4n��?�e�W̴�\�`�̹�g{t�*�~9ȿ}�9l},�Q��P������'skd�}�v_�w�!������{�.1�;�xhq��!��H�_��Ô�S�#+E/11�"���_n|o���|�S�e�<���6�`�gNy������a'�'���D� 7P���e�T��i������4�+?Y�s�Nu�ܞ7B���?L�P�|j�X%�c���eջ݈DX�9�4��T�`<���(0؋��F����o]�(3O��s�sm��y���%�>76~�v^$��c e����;@+��*���WC��\�a��B��s�e��Jٔ�<�4#g��-2ߏ=�3�Q�]��S� ��?��q?pY�qptS�ٔ��j��f��5��&����� ��5�~9����B@Zo��E�� �I�\-���(��{gA97gZz.�T��F��ː���v�\4�e�k#���/ J���}0m�� �Z���~ETX5ҩ�J~���7��ě�$0��'f���+�c e���6d��UNbO��=�bOyhٚ���QZSmW�����,��?6�L�����?����\`tD -,��Z�X=��NXlr�]\��y�w�]��"��PjU5�3���j6�^Ǐ�5�}R���l�6y�1qZ$~� Wv}�����d�%j�-�.�jq�E{B����))�̩�ݒg���N���H`'&�A�U����y�px�>R���}���t��DP"��I��;�:z0#��y�j՜���/��*�-'<�Jg��;�JЗ��nE�{O��C�P�]m����fF�����\����`� z��W����9�\Ѥ��ʒt|m�nF*��5Ӂ�6� ����9i��Ao��k�	^��=�6AP��YW=#&B�N�S�}�F�@b�p������N���/�rxiw[|���,6���]��3T�'�7��x�(EW4	8���nV����꣦M���O�0�˽~����HH�c_ �!7�H��[�nޕ�
��-^S�����4�������[�	6me4��y%6P�0et�n#�Si�(p�n��|AJ��x������}��$U@8z��2e��b�x��FL����jM<N<S�ʲU�Ɖ��- {nJ� Ņ�wX!6Fv|?B����2��z��z���ѢX��,���9��1�-�(l��lp�_�ռB"���~_�ou�b
ín��D��KJC�iHs��9����N9ܛ%S�9:W�LgmۋP�#嶵��E�:�h)��i��1I�����̂Y~�=$��?i�7WE����Q����A�&�'���vmcz��tJ����g����$�X�^��4�f�pC�/��O)�R���C��#���&`\<�ۯ� �=B�.\[�	����<J�Uy���#�Uog4p�Jq��Z�hU��b�vA�'tkRv6��Xkc��0'�8�������	c{n�E��h��h|��ߣ_�"����;��<�w]��x���,��1�����jW�?t�^$����e.���k�̓k�r�A����_��*	$�x"���4�9�M�<(>�n,6@�H�L��=���`�%��3Qf�� �5��w�����`�M�e�Г`{:B�}��G�cD�
&�9h����������.=����	x��&�$�G��a�^��R2��}��HADiSC!g̽��A ��;-��i�IҬ��);?��Q������}��L���y�U�ڭ5��HaN���%�_Ĭ̠�=�du�P{j3㨮��~Z�`���P4�k] Rb"-{h��AM]&��y%!����^8�o��Z:����1��6xҾգ*;\r����r�D���O����+��XԺ�nV������Ģ}Y`�w�@���)~+�d����=oy@Cw����N�XQ�[�x��a�n��3/u|�W.3��Ŷ`��3�De\\��!D�3o��4��tOTe�`Q�tی嗝�N��I���z`���4�:���볺����z%�Q���
Gh<��@ݣ@0���QF�q�L]祆t���ԭ��p��o�I�~S�����.�6��:N����Yt��قKe^NAԏ�6S�DY�3�8�
�8��t]����?U�#��,(F?�晝�(e������������r E���}N� ��4�D�Uҡ�Ӎ�%���ԑ	���XC����49aX����5nr����49�/ףs\��{$��Jl�����W�&�o@;������ճ�Q����b�${ؒ[!��4�X�w��h.� hlؐ��ㆨ�A˳T�8	x�/09������ȥIL�scC70KC�t���F�Ox�ʩ��^��4�\ɐ��tJd9�`�w�`�V�o5��P�kDN���:̊_�9\P�	�I��٩Άtw�>j`3X�P[�ˋ���:�qag��q>T��>h���D/�5�
�z"ݼN>�3Rqɞ�k?�-"��ы����������s��`1�����"�/�3
�~T����咧me0��OO���������Oߖ��/��إ-�X�G��@H���EW�Qj�:_`��0Fb�x�k���4�$�1c��/u_4����V'�>�?�5CUS٪tc�#�G�KuQp�Yh�}[��mM��jU�����p�	Vإgm�j�|2zޡfC������!J?4������f����g��59���9#>�{q�y%Y��!�[��ɟ[H�s
L�!��lKd��k��bsF_~�O(��<��𷣣�2��/�5�ͭ#�V��Q?i!	3v.�OiX(Fy��8�֊5c�����e�T�ĵ�`�g�}ψ��$gjH���s���"�J{�
������#�t�%�u����IC��w,�,drz�a�q�.V�?��� S�_���r��d�pB��KD�h�*f�����̡��;sn��p�EQ$e�@]����s��$)+W��P����8���̳�Cci7Yo�}	���vfw�yd��'t�m����*d.�:��N��iv/{����m��dwD�b=9�w��`8�%<D��5�Yc��J����dz-C�Y�������e:-:!�!�Ty�h�$Z������4o_�j�Z�G�m�FAN����T`b�3�کb���������f9��Wٱ7z}�1HvY���O5���~C[{
\a��_�����ʮ~��Ao�^��7��L:��EG�r����o�?1��ї4�����{�l<�8�P��iS������W�ijB���]���Č�rnҶ��	�<�a[�6��̈́�Hۍ�s�E~F�`�(1���lն��m��~;[�-��U;v�����w�#�9�ku��%�:>�w#=����5Ud1�⅑���)������0��a��:ە��X�E*zb����UwKg?��T�&�x`n�弨ei<��!Аj�w$�w������Z���N��m����l��=O�	���b���1�Tڮ)��H\"�	*��CGaޕN������9�vK!��޲���~X�C��C�9�\x���N�E|m w�w誽�jם��D疸*EY��6j@�]�3Z9~�}C��讀���Ɏ���SKO�G�tf83m,^H��V�3�ٵ"�Tb2	?tN�y@�4��q�˭
����a<�Y��[#��5{��hw�>��c�0�� ���If}�2�<er�ϔi������*��8�Z�{R
h��y�_k2�)'���g�R��rY�E����θ�Ɋ5J�*KTq�1_���M���9����:�A�k��a֑M�p�uvp�s�s�a�}.@Qտ���7P�Rg4��-���뉍G�ar+���O�&����|	'����(�f��_����KQ!J7.&���i�N��>�oV,G`x��f�p\�9eX'"�����s
��b?�� 3�YPv.��7�w���qV)K�k�@j�#b�6����w��iL���Ws�g�̱�8��3������k���>�o�=_E�D���
<�hD��&���	��mw�=斑��_qbd��|��9��O�����d�$�Ά$,��C<���K���\4� �����UM��s������| -2�GY���[e6GP�X��z!�v�Kj����	��&���RVx����k�$����[�R��d�����)RUv��g�d��Ԛ���v}��/ؐ�橣?eB~�D����S�@Sjƞ�Y_طf�'���y<�����q,�Gh�񕢠�^�*}VZ���+�2k�;�vI��"�}ɺg�z�vd��r��Je^���?/K7�w�v�I��ߏ^��f+(4�?���g$�J)���l�W_n9A4C���Y'i�e-�c�r�»6"�IC��fo5H~�礽�������j<-�M6x<i�D��zdK9��[�8�<+�2��O�)3����^�1#�9� ��k';p�jm:�Ȗ���|�1��!�r��: ���W�ik����<�7�c?!�W��RIbq�������/kj��"�"��g3�HY�6����/��.��x��)
"�)��3�A�}�L�O_�S�s��Z��~��O��q��f����@��Ь$�X��5k��ы�������j��d������{{0��I����;l�g��&��� }�]��Ķ<1�����ʥ=D�l��(�\� ȁ_�#Eyޘ��ωo�K����#ޚ8�-TJ6H����
:�h--J����ȣ�_~����2z�#�$n�Jm^�uO�3�g�1��į\���\�n���}�%l�ˠ��^ϾG
s�!�{�@�.:��a������5t1�Ψm�a1��u�l.�u�*и�KڐPk���Yv/S?;��3p��?�t��H��^�K���^��U)h��TRic7iZxASۂ=K�0,0K�8s���@5��@_���#���K����a����2q���<5:�=�H�XS���i���Y��2DҾۤ�*����A�'Z
�����a'7V����I�:���Ź4\�r���L�~������햌�2�� ~Ӑ�dZ		+��GD&/�Cݣ��ݼ7=W4��L��o�?���x��t��m5��\�L)e�(�cį���&��|�W��L�ʿ�K��'�J��*
.�b��ʁ_Ӌ-N�ڃ�1.�(I#�Q8���f���l��y�q�B�*o?��,6�u�6�3mk���Ԭ��q9�1V��t*}�Ǻ�K�y���W7XD�>��'��"q��F�N�G��;�\��W�XI�<D6��i�,�MrA��2+RX��Ƹ1LZ�l�' *d�� ��[H��ȁ�=����R�׶��៩T������Z�;1J�f_���¹@�7��j^SݦӺ��P�%%!J+�|���W�Y^{�%ȧǪ�����_����$�~����������3:L߾�����2i��M�6N$Y�>���`�Q�G�Y�Q��Ds��&�(��WKi���6Ha��Xci@���S��ݕ4�\	�RЀ���-��'��PL@�@ہ���> ���+ ��J
�L4&g�җX�Z�����B?2��5w�l��m0�<��A	���Rw��p3�K��'t������W$��*�[pyx<�s�RA��ۼT��-	�,��c"B�y^=���%;X���Dӯ ���(�αK���Bq�1?[�����ʨ��K����|_���<b�g٠UƎ�;CpdϢ'%G��W�L@qsZ�}.z��_˱4��R=����M0$)i[�Ԃ������N�� #�:������f����<�³��E��B�0�]�փ/��zVD«~ %[��TW�5�u;7�����(�Z�8��Q�6��3�G6m�����^���"'���)j�����l{d"��0
�M,!�n���K&�Nh�G�歭?��:S`u���_U��s��i���ϳ-�-�t���ky�^���PdW�3�©��޴p���N�jd 82U�D�]��̸�<��kcv��V��U��ΐ���[�?�l���<��?�}�?�`y)[�+n)��݂�s�`�%�����3��{r1�jݤ@��*Yσ��|���( Ď+�[◘j�oS>�!\�� �^��������?gh��W讚��D�(�
�7�`��ҝ��P��5@X��pn�co�r�����C��@Fg�O�>H,�r�h��p���/��Y�=8r�RЎ!�����'�{G��v{���O�#%6nq9�]�|U�&u�`з������,�W�;��>��-;��[��x�c=�)PQ.cZ��9�m�H`5K�+�����������+�$��0:��Z�I%^�m�0� X��������ȞF�O=��nY�=Hˌ��4�OJR��6�F��֊�-F[�I2�s���V#�n3��8D\e�p��P�^�d���+d��k$��.�l�U�o���*�?b�b"��{�A��j�r�-�x�3B�j�	y
�>�ÆL��i7�/�̏�wD,
�y���t�t�75-�4Q\������TOŦ~�:����\$��z~'8�+���/�)g֦�rL&�U2���$�k�X�p����+a�g����y >��X�q�3)XHo9�4�19��{y��G^Dj8�|WBd���ǥ��C �F�C9��j�b�ޝF�p.�h�>uks�����V��ުfu<]C�:�2��I2-������nDpqt!�y�v��3�6�е؂���z����,w�Y��� �?Ӫ� �a¥�A�1��4�ؘPt�9�q�������s۴%�ӤE}Y�.d���;hny_ &/�~A�N�d��`��5r�Ÿsn��g������yZԍ*L����?a�V�l�����h����]�
ȸ�)I�J6"|�X�G����Ng�Vn��q�o-0�0ݾ��A�P-Y�8��zE+�I�MP@-�h ��xY��ı	����@�j7N�
<�\�8�'�z=|���_�wF�|�S)4��F	��ص�:7�����*
��0;Vڢ��@0�tr(�^����,���۽�5�2����,����G<T�ԭ5������Ot{�i��_|�|(��`��<9�fӒ{����\�i�i8�������<2�cV�AQ�A�s�����Ɇ�������r�|뛀�qV��q�",]$��n��HQ���)�t����n�R6���u��iZ��_��A��b1qV��6<��c��,b6�Q0���R[n������<�XY�M�F�G�3v��_��gz"�!�c˼�:�qv�-v�g|~�RN��b�5��G�͉B��i���4Rމ�<9W$�վ�wz�WV�~6�mq<��UL��	c 0w���a��?FYrϕ��l~��t*H�3��y��0�WEʟ���{�֋,�`H*TyO���Խ<I�x��jO'�j�)l~)N\H�կ�g����\s�����E�'-g,�u�����Ǿ��n~$��Ƥk6iLT_*��`��m�{�!��@��?CH<�\��U���3��O���˫}\pg���eHN��.�QN�� B*�#ĭO�Kq�,�#Ք�%�@[��[܍n���A�&r�uk��2�=2?�s=���t��-K-�����S@�(kO��6��sl��d��(h�����+��)��(j�0Wmx�+C�������:.bp{�X������@md�.����`����'�x�@`�:å��Yl�� �����PL�g�b��mDM*nk���Y�ҙob�c���&����v񙖕�\K�H�&��6�3�Z���rj�#��<�DOT�s�x�� ��-,F��&L.}彉�	�C*���Z��|Lɩ�L�ӋT�9L/���_?�2�j;���U�-�N!��Y��U� V�� BĩE� ��}���ب?���6��(vh��Á��g�Ա+ -��mZ�Bmq�'����e��p��j��%@�7?e0뿶X�Ӌ���k2��֢6����.�IWZ�m�����Dsx����l+Z�(�9��v��<�Fp�Ø�E9�(4���)�%�nk�i��ma��<u5�.���m/e��1�ND���G."�h�-�-�$���_o�Z&Moe��>e��P�^�?�ԝa���fQ\=$�$:n>y�8��VRc��8��,�o4�<i�����]���@�n��	k:R/�B0�r���&��߈��O���a�i$�h��φ���<��z��D�ϰ��4�p/�R���zo.�*�*` ������T%ZQ�+�+�o���zu��r����~�F�g�0�2���474|V�^:x*�! �$O"'<���F�'�M܁n�Dn{���RY�Z��F��O�:�>�Ϻu��W���R���Gxs��;>�����px\{�9uU,[�V��<�9�v���bl����G6��qO$��?�p�H�m���B������P��L��v�A�j)t c)��D�z��r²tEGE
!ˁ�Lni%S����|�D>;�.�ۀ�:�L���d���$�������U��p#<p���3��K׌[=#P>/j+>�mN���d�ԻΫ�z!8�����V�S>��l�EZJwy�l�	���|<��I}8�~��өJ��]k��b1�}���{��X'O�*@����{U>1�TF��ܤ��_<�u���BX�>>�"`r����,��gL�t���ʷ3����q��,�:��`O'sJ���N��� J����O*)|�C��A<����N��8�9����5��9�u��Ē���O@���1���"�C�~)�k�P͆�(��������J郠�8���!��
B�'K[�b#��
��͞k��D>LJ$��dU;x�����W�CҦCW�r6'�w�&9�=�(]v=�zZ���ƪ�1Q�j�����Я��=C2�}�N�3w��fCa7<K<D��}�YML���?N���
��U�R��fG����#c��c\RԴ���NUH�A��!Ur�;�&���t�Җ�_�� Wغ��G�̋��N��2n�] "�V��0������9����1�)�6��7)Bxdܗ%_��{c���2Af�Ľ��{Jt��A@4�%8�0��<�:��\�H��q�n+�V��BN���w����3"9�)�nO�G��ՕՙJ���kjP�� ;�A�âCn�FU^�"��
���ѫӄ�`,�<<�r��� �V�0�o7��ƙ}�3�wKG��@�a�]4{@BT��U��v�Tҕ����pY��7F.�qX�%��:9ռ2�F��˂�a�݊4��7슟љ|��g��*����˓`�PvBd�'&*��
�����Ҧ#��&����I����4ĉ�j���ص:�-��5+#ф���1��V���)�	Z�45"�T�l������݉a~������OZ���t��\�+o���V"�����	�\mT�!%)`h�*�1���/7���8���kT�5<����=Z%5|�K�BK���~]|ݸa���Qg"E�0h4�J�6�NV��9���Z��\���_Q�ޜ��f?v�kni)&��}l;I�,s*M���b�����V�������[�5?un��{�gW���f���q�D���,f��T�԰_�X� �^B{CW�\_���sة��)B
A)��t�NP�թ��Sq8�4*�s��.�Q^J#"���5�t�#Ƨ������v(F�d�����:Uw�,̇/J�\�4% �b&�EUH�t���gEHz���dl�6��Ͻ�d�c���-��^�~d�4�^���7ƚ��������Q'd,:�������t��0��F7�=��h��*c��}�8�B���l7���D�VuKK�6�<�<~�>s�Wr)�Q��b�K��zO�[�X�����Q����gg�/�}���2�ZN6��/U@+1%0��� U5ă�_�wZ����C��b�&�*��t�1k?��������ĳi��A��J�ެ�rn���Lw���5�B�+�n8O��J.9b����A��N�߰�v��*�;	�E���:�t���a�,Ӻ��	3����E-^�oJ+�c�]���4<�`b�W��٪b����T`B����#��q�!i��&6/�x�]��{�>��ͅ���89Qx����~�������P��r���:h�Y�l�k.��[����9>�4�'ֲ�O���״��E���ę�n9��-Cop5�T��B�L��[��|w����)�9B������2 l�sg3�i�o���2������1��p�����*�T�(��x#���ƒ�X�ds0.�f�Pȗ��@-��<g^Eپ�PVU`�ma�+K^yJ@�
s_�i�M�T&�����Qm�MC�k�C�x�/ݷ���a�UE�t�`�r�N��Uv~��LxR��$�şX���4������ԙ�Q�4cF����?�ø�c��~]�R�-'Fʑ�0%���f�Y*ը��1x�&�q��X��=5���ӌ bT>�(�ib#��Q���_�>h�-Ӆ���	�x��g��B��8�����F���h}֘�Q���ќ��ɖ3��:��~��]8;\�����l�o�$�_1��w�<f�l��O���I�/ ��:�"��xZ�)�/��9����ŭ�-�л��q[
��9Z��� ��aZX [?�ݟ�C���C�%��� ���I���P8{��&��ί�h�=��b��{��G���d�{�3������i�?�.!���+|kB�٥��X��v}����#�`v�\���3���D9�|�"���-�'�a�!�*H���<�	���[�zAUpԬ���SbG5w�5947Q ��SKs�|��7��a]?��M�g�M�n�<ӷ�*�J�����oh$�>rp7O�"Nb[7L��qe��N��Ȃ��}��\(�-�iG�9�Xu��80�|x�:ˣQ��� ����v���4Y���;������d#e����3$~�݂�&!�r(�k-W6���gK
���¸\��҆(3�灨�������+7�,ǆ�1.��,�f]�?(�T�<�P���Ww)7�f�ts����x��'��זB(^[�F���wL��6Bg�rB��'ڤ�@bb��df�Ťg��r��u�r�j/ٷ�@��AC�2U1�=,�e��AU!��M\�^���#�5���p�*?�\ E�����.�D%&^�h=��99�B�)���t��DH�us���U�4d"'op{�/����t;T�)P��O�gşb #b���_��<��L)�+2S�s���ۺ��r.C�N�UG�2gkn(~���6����	Z	�Н��#��Y�������v���b�s���ڏJ,��v�b�"�ﯹ� ����E�?��]��:�%I����PK����F�j"��X��/�m$��߬�*��T|�#��
����a��m���=�Yd-�����s����g.rʘ�nL��Z��W^��&*��b�@���N��2��T!X�G�ю�Gk�|�Ɏ�:�d�s���N�_v���$ "Ɠq�(k�)
K��2W�Ҝ���B��a���F���~���ӌ o2���,�bXX�P�D�	tゅY��'��[��7������ 	d2�v�тj��Tq����T�J�Ϻ�F���L����f^\��]S�:�oE����!�Y��tv��6>ɴ��:�4�Փ�qT�֌m'	����O��Q�����h~�&@w)��6U�O���su�D]�e�����gF4^�N���7�β=+*\�$� l���1��!.��5�:;%�jB-I�P"������|�{vf1F��B��m}/o�NH�����:�gH�=�Wq�~q:�z���W����D��>�΀�20���ߧ���b�N rQ��#uY$"�+��Ņ,��b����y�lk��tt���wh�i{>���!����-��b�N` ,� �c�h=$!����ī~łX����j���d���(k�I��5��i�E��^��23�P�W���f`%w�ެ��u�`��L��tv�&�@�:q��3��z�h(�ᨊ+�{��/��Q�~�S�a���O/$����s�*�:��Qo�T�k�0�/�r��Բ��[���FK�H� ����xC�i�������y5�\h:h��?e��fg�DJ̀�Q>����	�M�]�����wL�9Ba߲������y����5P�rr��׍�#��@D�@��V�דh5�s
�d��S�4�ѐx!qܐ��zd�E���9���^k�"��� ���V���y�W�k���28��2L<�a��.D�������|dZ ;�-#-�'D�'u�������.ƙ���>N�._i��HFu�� Qִ���瓢�Q��
 ����F}�|��.?���J~�7<ٓ��U�h0h�c�w��L�R�(�l]���8h@v�)��Sk����Y��d�c�oJW�P�����4Ԭo����Yw��
�ܸ����^��� �����I��#�&���n��y����~�ð�-Ѫ��HZ����)��ܶ��'U����w��^�,����o ^��Kй� Ƭ��[E��cpSQ�\K(v��+�d�W�Bi��b%���U�ƿ����h�� E��,
=ܐKάP�*�`��C�������9!�`�{�t���B�'�/��:'#���w��}T+�=���c���S�mھ)�{��Gl��_N%sM�9��)3࣬'zB������bO1"$8!�5���*S���ȉb�I�S�~{��t\�i�<�N�2W/.�<���C�����:lh�У�,�r�aC�¡杙�>�� ��B��w��#��7b�&k5����[2W��˜굾q�x������G�dbo�<jO��Gg�۬KL��Y=Y�-��(�>f3�O���GYsx���Mw����g�(�=u3:{�팭z�P�_�5��X�~ۥ ���+V.;��(h�`�3OZPN6�[��9f��w?�-����,:ڹ��%v��iMa�t�K��X�������\������Jb��*��߼{
��C����Γ�1>j�׿�譋�ͩ�Q?�N�g/d=���u1"�p�OD=6Z#|A0��,!/:K��ʁ�k���w
gLz��X/�ӫ%f��Z��4;��o��*ЏX����;Pp�ts�������0d/�NG��@�cKmd�_� * KP	�~���31�iZ�	U�b�D��.�{&b&�A����]A�������\�hN��ݹzz�㶵�#nؠ���$~�)C>��ݹ��.O!�.���O�+p�"�%>�Z��Яb�d�^#���ܖlo缐l��'/�~	n�%��*Z�$����qې��(����Q�K�e�GC2�y�L�w�b��ˌ�#cQ��puC<�>�O�<�9�m�:
�չ�FDGZ�Y~:�������U�zG�O2���T��w�ߑ'���y� G�����yq�oX��y�i⤞@����͎\�����B��@�[�%�l�ŋ�q}��@TAP��v�	N��Q���������I ��1�.�Bh��ƞ���|�5*������Vm�k=2�v9��s��ݻr��8L��o�|�v�@���,�~���ߴ��kh�(e���̲:�g;�0�M��-�2a&g��@��ɬt��j��`D � v�m7}h�\3�l̹���QH���Pt��Ap~A���ϒ����T@��/����0�U��O�)`5�uǫ��ecnwqg��������sn0�w�S�1����'�7؎*ޕ���-xZ�Q�\ƛ�c��d�4��d���)�%w!�F:7)Ӆ�7MQ4�~�T��t��aIo	P�W� v��<���&B�o�y�;�m��0�RFT�5�	�@�U;��Qh~�6������+���m� �8���}c�ز0�p)	�^���<Ǣ��*˹� �P�S�Q���+�. z~}@���HT�˖p��!���`���D=S��n��_�����N�<�0F����ܟ6'(c̙��a`���>B�؄o�ëw��gR_D^�P���� =�����$m��#`0�+i���j��I�򔋁.W���q6S�3L8e��);1�v��Fd@������L��t���hFW�J*�t��n6��p��<޺�l.���O���`D��_��t*�pcv�*�$��б� ��>�Gv�o�7�w��I�B+-P����ݍԍH2�Q!?���|!4l(����P��>�� B�&^����i�n���20w
o��CzN�S�'Z�ƺ��+�L���� 3n�V1�gtl�q���~���1+GL�۔Q�Z=B������Ԛ�X&���4F�n��!�r��w��N_4���v�߂29n�|����&�*L�:	\j�}ua���p��*= �zĈ��/
���<?%�O��}�Jd�:G�4()�o�9V�D�Ƹ��c�3����D���h�����2��S��'�����i�@�l�֍��t��zwz��4g����fT�>��w���CLd��������l,���׬/��1n����@N�$�8���i��=�C
t͵+���.�Tn<}Zk�c����fhl�w�Rݽ)x���O�-�F �H1���*��F�S���"#��ޜp�p�/2�B���C��9K7.8��]�X����<J򼎢�K���������r[�N��}�[oU��K�e]S	x�O����|��h�S|��>�h�,�r2�nL��:�u��ۻ��X����x�)�uv�\:U��e�dt,�ǀ����T�� �T�v�����<q���\��S ��9���HA���>���କT��i8*�C���P!Q:�Wa��e�/��2P�Jg��*;<4�=T�c"=���w���U�zC���x5�z�GޙWM��?hz��}X{ϖ�ms?�J���M��"*Z>c6�^d-�_�^>���.���#Ӽd
4@;���찓�3-7�2yw?j��Y{���ȥj͒L[�3%�|0�~��[A9y\����z��I�o��v��O~˺(�I�S�nf�i��>0k�4.��hK�Y�l�_�ަ`��崠A!ݣFD���WC2��2t��o�/'S,&t:$F���� ��|���˳��Il�� ��n����,"K�b"�w�z�����Ҋ�G*�$)/��,�?�9��7 ��>� ݯ�_۲�y=��L���]��VX��W߉z{?�Cy��*c&�sS0�=>~��5(KK�T+^s������B۠��n��cP�	�*E �ƭ���bTŖ�5<�՜Vǹσ����o'��+
�����R��e�K
�
ھ@5���&�J��$��<s�+k��װ��(���֩�JL��HU}��)U!�¼(�.�#O�A�*:�r��T�	��2�O��3#��-�H񭵺��e�)b$i���A�-�X㦲�$�!kJ �Y�1�^�l��ڈ�ֈ�[P�z��E����Ϙ�>|���ӯ蕁�d8��ОvM��8"�KƟ9k�����}�(�sK"_��iw��/^�����rs)�x����-�~6��䡸o��	~��k����>	�������t<g�y�,}-���-"�E��g��Ѷ�L���t�c���9�v���U5����r�d{0��)�3�SN��|���x?w���4RLZ��2ɦ���f鮾�ORZ��+�����7~���W*I���Wl����h������'m�"�������5|K�$��]}�f>uxa7��g�'��Fq�A�R���J�N��֫#��}N #Й���g�����p�vq$.���t��wc�F��B#�8��O�˱�>?�w��ظ����ݕQه��v�dߖﺢ�lF��R1d����ayk.���g٣ �SM�v�]���ruזq�(d�6��am�~�t�\��O�I���Z�up�贔,ߣS�Y�$�SҕW6pv��V�! V]&{i����`kMC����8y�Oxϋn>k�f����]��|����ww�c}�6���/x�Kc��)�}y޾��J`+#�nS���C�BQS�X�����#�9�3󻼇���3����`��9����x�?ҏn���v�Mvh����=��h��ʷ��/kg�o��aI�h7*�W�x�^�]�ZZ����͊1�2s�0���l�)ʡV�����.'k�n��4s�E��)�i�ǹR�J�Ҩ2��X���p8{r	�zo���:6I�=doM�%��q�_6�g��,J�\�3j����FZ����`+1��ÓB�L`T���}���g/ks�ɤ��R���13Y�|��-Hx�&H��(�*�l�y񭞺/��.�	��vǯ��a��u���Ȇ ���6=L2�I�	#���Q�PB_Sw�`�iV0U�u&� ��S�<>�k!��[x��%3�Y�~u���Fy5GUJ
�Lr°��Γթ����ObMn�j�@O	�Bl�(�=���lу8�ll-��fE�ϫ��F���G
�'o&���r���Ѝ;��
J+�Θě��peel!�U5^x|�(� ns�G:�*U�z(ґ�����R�v(zN[ݿ�C���J�g=Հ��eM�?AT�P�iQD�AИ�sϡ�5n�E4X�J�)�ƅt�����%��o2Α��gڟdm�_�#w�Fpȩ�T\�Z~�j-eO�n�-h��¹��㸹]���V2$�CA8=(�+i��B���W�^3HS��D*~�<��]��\���)���C�3�eZ�Y/˘Y���r�np��1�z��
?���!�cK^j��h��6Ƌϯ�s������W�^�E�L�&	�O�Y#�l�FgN �!d�~��*�{猓��:]䀆�9OD����-"������w�/�"E��N��8%>�K�N	~ML�}�|��:�1��������"�n��R�4�c'r�!*x���a���+ŢmB�t愂�.L��bY[��W/pz�)Ü��gI�-�>B2�����L���H����-�2���Ȥ�Ë�m�>$q�g�
�f����	�V�[���[3�rj;��|�}}'H�<\�Z��@l�����aTORV %X�:%j������'�w�]�uX�1*�X�R�٫45'��L�a����#�z�@C�Ҿ�8��q�v���<��t�+�����	2{(G�nVv��zhe�@�ïl�&��/��ǒ
�af!����Xu�����+%�)�A. �6Ԧ��b� ��z�*�?�=��s��F��//�}��m�aI���:I�8��
݊zC����*ƵT�|�Bs^zR+��%�D��𔢪�h>��4*jK;�-��
��YC �{i	:K�N��_�k,]�'�"���{�HK��5,���x��-7��y'/r�!�|� �<���Um�Yӻ���I<>}�
gW������dʫ/[�3��j ���u�bJ��MM=YN��0��?���r�����t�qɎ@��g�2s]�6������l��.wg]�M����%��B]����ȿ9`/)��2�k�6�Y������u#�<���U2���q����C�FY�;�g�\)-����	� =)��ƶ�|:P%�έq�q���=�.�3�l/�SD�e���W��?�cw?��;2��^�?5;�@V��Y?��&%��5���n'�ǿK�w�:$�CjI!=K�Y�6zE�QF�>Ż}
�t�A�G�������(~�ӷ�B������L3������^�l�O��j6�
�O�Ya/dڮ�;��/�7�'�Ӆ��f��<ը��k�M��p�~��7�!i�{��#�Iip�)�ЉL]=�Z��o�k�H����py~�_nft渲'~� ��j0"���D��HAﲝML��%�q�2h!La�R��<���{��4	��|~ �┩q�?��ܖ~p'��Ąl�<;�v� _�ň�~��h����Nt�a���������[p ���#�l�ⱂ��kﰗ8eӿܠ?�Y��BUmp��'01;G��,���8H�Z;F9S�YC�� ��q�:֡�Cx�������P�M��O�z/��H�/y�&�8��2�C�O�!�2֝Ӆ��M�M �w��Q�5�h6��e_>�uj�����]���t�F���y���z�<o_���@<Q��ßw�fae������f�G�&�O娍Y����+f��� T�`5�P��XBO��#i�n���Put��x�'���@�R���y4HB�68ri\��Ӳ5�S�Г�n�Q�,�O'��O��qP#�N�$����r�ɶk�B߁ �~��@��,��rlc�U�T[�p4v	d�כ�#�.�� ��Dw2 �%�LX��3���*��*(�r&��{�ڂ%�U/Zy����(a�;D��Y.ot�X 6n5g�{�)�]������g�<R'�jLZ$�7�P��Ԉ�D�t�0g1�`�/#g?���@���2-��%�:<��4�+c����2a��_�eYZ���4�� W�����:��a�Ŏ��b.���s�ӽ����R��B�!�����E�qo��"I�؝H�� �KS�`�E'i$z6�+���� �[2O��Q~��ꈳ�;yFk��)}��4H�����B����e�mlYOC1ʋ�A��V��\,[Q[]_�7mЛ�p��QS�Ơ!AZE�~���G�a\���KQ4B3���+7ȥ<O.GB��48��)��/��� E<���
��H��9��@[Bt�_
y@���ڍ�l?��t
�����g�g��W��M����O�-9�'ht'�2\�E�F�{�SЀ4���S�O�h�^\ I��
�^����ޤh��*Q��Пd�/�슞Tؙi'��FO���i�Ŗ\�ܪ\"R�#��F
0UQ�Ia�,�0����� BN��K�DS,��{CzV�r��0�6��MEV��2f56�>��+/�%���9�I�T����V� #҄Abc��R>�?'ō���;�^����Ŭ6^
.�y�w�O`�c/�JjZ%=|�n���t1Zp����lUY�*���}ؒ�y܄ROx[�u�M9漣��L��qp��������Qcm���A���#T�l�lOu^������6�S���_vbb�l���k�v��(�3�-'�GZ�w�y����AF���h�G�n5��xS���s�CƜ!�����%�M����Y�I���/�.���ۚƀ�р �t���Kѳ�d��qLI��J����^7���U�����t)�9�݄ώ��-��ڈ,����iy��RA��q];���:�h�H�tꎡ��~DMD�-�	X�Wk�t4��)���`>��B�6�\w������ k9�õ�ug����J�e���B.D���+�?}Oa���F�\��Г�~� ��)�KGl0|P�s���5�\��Q�r�����}q��_�����ɌY�+H7;8L�O6�1?L�T�$��JK�}vAG���M���X�L5?�_���us1��<��Ve���m}��s3]� я�\\b^qES���Ejn\Rs�D��N$�]ſ��|� o�_�P���5���������3ws��b��ԇ�x��]���I��d<��܎�F������+�]�[�݄P#��~U'���g=�}�o���ao̓����2��VA$f&����*bUnV�̨�z�6yqF��w��?|$tK�(�$Za���|�v��xYx�4`����f�K7��oV�:����L���k��Oi�4�Dd�8����%��>�/�*2?eN��Mjq�v�)����`q }}!$K�^�����
B�x�Ԛz����r`��0�R4]���^����J9�ޠ�E�l���@�q �~�1̗aw~�1/J�"0*��]՛��.<�*%J��߱��.
2�a�1�9Y�Wŋ�t�n�E?'L4�LOb�T=��~�l�ȞA!6�u~���́G��z��X��D�N�)ɟ(e�&�;��� �" K*H�vGٞ�{`�R#���rA��h
��8�\����9��������/�;)o*?l��t��P�+�3��Q�6�z��
�+"mH~I<~�;;9���I_Q��Q�'w!��ʿ|������5i��j7d� SH�@�W	��WzP�K/�mJ3�k��X�E#S�s}l�Ɯ�Zp3���ƴ�� F_o�f�}���\L��3�6Z���N��F1�z� ��^����,��:��`�	Y#�Qq�|�u����2Vc�x�D{��K�v�.C��b�f"H�������ea<\���ӻ�l���hx�<�t���"�0�	`)?��Y���m���S$q9v��tD��{E�Q���X�s6IJM6J&.}�f����ā��Ou���h�Ʉ�Bk�e���[3Ez�Yd�Rz\pY�:չq{%YdSf�.�Q��yђ�i�J{"�|���&*���["�DͼXe��lo�=����kQ�Otx/ﶠ�X��~��c��P",���Y�s��xm�O��ë���=��l=#��*L �g*��^)�J�~�Qہ�(���K�یe�x���$/̸�F�S�F����B�#��ܾ$�[�㯤򛋆��^�6�-�v���d�j���w(�6U��ˠ� ��J��-�T� �஄��ɺ���FR��m�<�0���S�Zs�FM5a���2"� Z��F�r��_���{(O�����#�@��l��WMV����ki���ͷ�/�6��B��b��Fq�]��#�j��m�Y:�3x�	w�By1ޟe��Zh��nY1m�(`�~��'/�U �fNPG�#89���R� <� �Fg��و�)ǕF�˄T? �Tߺ�Ap(!�>�F��5��L�&q���>o��.#�aa��J8�&�9��p�j3�?5���aЪ�EZ�B���6�_nc-3���z�~aM�%��S�x\o���r����;�#�s��Q,�l뤈���3<��H�;���~�,�כǸ�/�9 X������$�z$�|����-q��������J!H�Ul�����]�\�Z
�'UdF5l�&���%b5����6��]�� �OȂ�T��͔)���h��0�L����`6��%\���Ki3����|N�9������B�G2; ���J��i� b�������hgA4+��ཧ=��}
��{9�W����~����H����fjx蜳����T؈���Y�a.I����q���D�>�hF�Nx�W1���&׬�_e\�D;zR�t�̄�aUK�5�� ����P��u�1��T��Q@�� ��v�- ��/�n��|Y�_�;�,B��E�0`z}P!�\$㧋wSF���rC�R![�R����eO�L���
�Y�G~�Ǯ�<��-���DP��-��&%�h��Z���d���:��oɡ	�-���Kgv���n�� (m0
�Η��	G�k�)��p���Zz��lf#��{����C:U��oC���i��!]G��r��֊q5m�&���d �5�I��(����Z��s�
u��U(O���VJ�ź����cr{/��Jxw��s$�l.r��^���a��RTp|�dc�xb�͕�k����S�������ܨ���f��%y8v߲vO���	���a0�K �Ep!@ׇ������������m��� p�}L>�F�~6s;�u���M��
8�d�<F�i��M�)UӸLg�a�2qQd�5B�ϋ�!s�M3"$���/�)_`�c��/��-��L����	��= �z�\fj�:�GTWȊ�ф��m�D4��n�yk�1�%ta�a~�*�i���U&��7�e�F����'��M6�8j^��AHn��G��?u{k]s���=�5�����E���MO��`w�D��Z��J>#v�Fn�.l{���AX��ɴ���t  |��3$'�d�jQ�k1�Fa�|�O���UdH�{���P���� F�xb�}I�?[�J�υh��49�\���?b���,�\�k��^��)T1\Pz���G2��d�X�yИu�/Z��{�m��c��e�M��S�~���`5��O�קb��,֮3�:l+iGG��\�Q���!��-���H���hwxc��ko�(l�$,��W,$�׆)�:	�����y�Oe��8/x ��N�}���fw�蕮<f�e��O���΃*�ShV�>$] �t�iIs܍M\Uh 1��ɐb�5/��jh����!.q`��W����ot��;�6�L}��1	l�kM�lv=��^����O��U��ſ��wl�8�[��m��R���Ѹ��2r�&/@�����W/^��k��!t�~Og��w��{6��˅~L��?�X���x��N� �,T�Шo_^�J7)&��OW�S?]PXűu��X+��V�Vf ����t�m�C��N���n��x���Ѳ���2*�|�οI*L���*+,� '�5xRA��d	��
�7�<���"�����-�0�v{����bK����؝����D��
�{�����d��W�?$�T5�_�v��;*�K�Pu��f�
Zq�䯿���a��|�!3�R���@�fpy�8�M&۞���9�EY �7����M{߁�>���V�OE^��湊��ѺV]\u	�}tA9� ;R�5�Fƙ����k3rij}��!;��'�R��` ���-q P$?`��`h����C���Y�����H2ى�+��S�hof��%��0d2��5��F�O""�'Ӡ�]�P�p���F���+�*�<�m`�V� R��RB'�[��I�-��T��\�z "�iR���)��In�J����|r��-�[1k��Sm�C�:���ç�Ve���c�� �o$0�A*v}j���K]�3����r&��O�ٰ���3T��0y���*�b����v-�>���� �2�{B��|i�
�L�;�msU�)cƟ�	eW��ķs����+Q:4�����i.��ڶS3�E�����$�`G�E�pL��P��>*�z�M���Y�D�Y���I�aӕ�����FY��͞��ED�8�|�?Zg��q�v�W���!�A������w��}x}�ȍb������`_�H�,�6�q�c��.��X���y���������{���P��a�&�1$4�P��E�U�X51PE�^���+�(�Qʣ����:l8����g�D�}L����W�d��S0R�W5y�����f(��w�g���ڠ-�]`����Kș���`7��"�	y_� �g��D�/�
�UΝW���/3 �X�w~*֝������BGK��c�9y���w� ���o���«B*���_�p�Q����-q��Ɓ�τ�9��
z�-O�k��Z��N�T�C�W�����?)`��x�c����}��RhċGp�Ez����!��Y�Np?�~�/�\sr;!p�M%��� ̦ޣ5�ɧ�֫P���޹�[������3�$-�z����o6>&�7��ӽWv�l�c������m:Ɏ2����V�+:�AF١TS<�]���8I�C#X�<���!Ʀf�W~������� ��4 �0�&�2�)�`���o�%��z7�ޤo뜈��������%o�R(���[�~;y̅����'�>��M�y}���3����.�@��[������
.]rH!��c�,�a=���b��\���%����7[Y���EC����k�^�)D�Q^稶�Q�㴀S ��@A|��W�ϵ迢֝�����6Q��'fx�N�b�N8͝~��o2��FX���~�
����xSd�gy��LL��?���R�W� '���R������my��.Y~{=���c�F��
m�����FxwҭF���;��}����9��������~���3[{��I���l�ru�r��S->t����1w&<b����W�a�E�j�n���џ8�r]���Ʒ9�	�e�nP��>����fL��*5P�Z.��.g=�7�?!�z���~�!���-v,��`Sp-���`r��AbA��
��R�u�<w�Y{�N@�af�c��L Z�Y����6	�����b����W�R�C����u�E�M.Tn��r�x��7�W�S$R����w�����7�6���	d�E��60A�Cd1p#XY���M����~�'"롊̥Z�>�p���aX����Z�����2�^�I�� -b�]|O��Ǡ��"�`�7xz�G�
��y	�NA��@)�~���u)���PA��+'j�y:���^�RG�� ��fk���6U}c}cxAVs��֮_�����1}���&��YdܫeI ���n�'|��Ts�۲S��o�󠕴��O�b:�����{��?�)L�%�����t�t��1anz)e�� /-���k��u ���s!C� ����� �s
��$R�<���wsD��JsZ1 �$�/g�;|s�U�o"����{�|�U��DK��N>��d�<�58��9�c>@��~I�>봄�E����W$�"�u�"7z��C�\8]v+�"�޷g�=�fO�sH� ������9]��ܪ�N����ҿ�.�u���"٪�ޓ֟񅣪!�w����K�G� «D���LE|n��̷CF�� L��ջ���@��/��nkG^] ��7��'�3�W��T����� ����J�ӹ�d�Ǎ<R�l�d})�c ?q߸o44��� �?�XL��s�U�����Ɋ��z�4G	3����e2� {Eg�W� �?o.;��$7u�u��f&w1K��^��E�"��f"4;�	&j_����rU�������~.IOb� ��iv�_F�����D��O�PLXx�|�V��XV��4G==T������c3���V�`�y���V�QCC�����-�j/�BJ,��i�A��zE�v�W�Kg�`Ov8�0�%k�zએc�(��eP�2D����H)D��D�ϾB��W��Ⱦ�rj��k�c�b��R`-�(��x;�I���������
Weyw�PTt�����y�h/���B"'�#-'.n�q��1^�
k'�Șd�1�����8�Ձ���&�\}��VvMv!m�����t��a��фK��^�g~�FZ�ܵ ��f%PL3kkp�;��*X�����u?�`�l���=+B�4�W��8�cS�O��C��#U�	���n�����8P�Q@E���#ĝ�~
"�a��U���h�ay"emY���<+;7���k,j�)|���U%���=��;�I�G�������f��*6J"�G�:.�멹�dS���ޙ1MZ�.ǔ�Sc�LLWhW��D�J7�!;
���`���;�e���?���8��k��N����rH��zO.��0��Y	��H�A���ݙ�;���,�����^!�6�b6��(�_G剾*��`Ӳ���{�>'�2���lG]	��29�!r �-�mU�b������<��[��<���)D��~_k1��S �~�碨^)��X-���>)o]u��c�#�
���}�n� *����\WxG!^�z\�_�9Lr��9��uB�) �-���-�|R�uvt��7�\s?u�%�q����#���C�Z�Vg}&�88S}[�;�+q��5�u���?���kȗ�>�w��v'�(v= J�Y�ZJ�� W�n��P� � �+ѱE}�M�6d�뺵��I��
�ԯDd����-����>�'�Zv��)�4���vǈ�cO�0��>d�h��J����yu?�,��8���A)~����h���O�X���)�V4��!�*�uAr���B!D��	���O�D�ʴ��l��FT6Q��t05WV=���_�᥉�'����cƷn��/��l<�����S\EA�p��WA�߶mؕ��ִOF�+����SO��u�%Cc�ߩi�s�ώ�*��v�WSVeRIL�V��`���5e9w��V���-��P}�n�ґ�����XN��u���p��.^�d�����Ď�X��~ϙ��i��守Ǚ���=��)�%m!:?����G���S�h���.�$f��p�J�וHٱ�b�z�yFcuQ<���^�xe*�,�%��^�(�w��`K�����d�nIO�U���~ϱZ2@��Nf���k�(l�rz��S.�^ �uW�=#3RDXo��Ur�n�=��W?�{`��j(��n%���?F�lZ�������`�n�]L*}�^����t���4+ݼ������cSD��H�6�~A,���k�q������òD����m�ow�|�n�Z��yNŖQM�O���TR݀����o����v�A��6�[�*�
��z�eq�(�8���6u��g����%Oz��r1�哱�qp�Ɵ�܏��Ґ�:*&f�5K�;�^w����k ��
GԳ��<����`�D�A]��Y�w[��sF���|��%!��P��齏='zW�]�p���~�Vox��C��j9����]O���J(��m��2r���m�ZE3bR?O����(�}�����_�S�w���e��P��eУ�&��	i��z��=P�c:��Q
fi�J��J��X�Qy�9��:�/�I̺����z*��0�A�"�&.7W��;����t�ِ�n�k�P0���_����Fa��ӣ	� !���5`�����m��6L�u@6/l#��4�u�v��[�6"<)u�d6�%���b��ь�+(�������Չ��G�vYp��_�>P�:�+|*G�N�&%���~��m6�C$z[�[vՎ{#�����g������3&F]�m!<�ʿn���n�G)�ضl�� 4����&�K�`Ev�E=��8C�W�7�����k�L{����Nh8��X�ZO-����R���\�"�~	���'�ՠa�G���� N��i�V��?	��S�G��㠃�Uȯ;j�ړ7˶����7��T�S���K�T4��#��
iD�i�gvR�UPs��HBw��K%�1	�%9r5� ;�o\���tr�H�jv����i����2�UP�5��#Y�Df�13o�F�}�P߼��YVd���d���,Q��L=�6����"�����"��Z�MloBvAS��Q���1ZR`��7>Ҟm�x^������D�4��!*���!�HaO4�ED�23�N��Ϊ(C3�>���F0��Kb���%:?5�0<�Cj�i��\)6g||n��<��6|X������k"��w�\�f-+�bNrk�sSJC��T7�����q�&�\�y����D�{��r��\i�R�R#s^8�T1nY�2�f�(e�-!L�����������"w)��{��� �L;{^I���0ѹ9������X<B����:���@���� �F$I���l��7�}<�³^��%Y��<��t�RM �hI��( ���_}rYD;"�C��	�����I��,�?��M����_U�G�K*@��y3���}
�7'�B�T�`z�@�[ռ�Z�Q^^)��$}X?#ю���p
'n�	���[��Q�]���*|
,�~ ��O��z9]�]��r�/�Ws<T��&�y��4�bÕ�#�w���%/,� �vn�ټ��l�f�2Xĳ�5�Y`kL�ǁ�@��k-\��c]P�r��q�n��H@_��"P�~VF�Vk`�+�d	�4瞄tEl�Ym�v:�u}h%s�I��G\ILӤ�*��1��OԛSC�9�D�j���Ƌg*�k֥��Q�q��zJLg5�f�'��v���i������/{ӵ��_�<��y�$� �Na�"�s�
l���J2�)
��q��;Ғ��遱���
,�2� 8e"�TI<�����ƚ�C�HBq�ŕ�fp��P�;�^�� �+��tfC�͸%��B��MPvpZ�a��+~Kp�\� }ޤʈ��}�{�W�g6D-͒uO�q���nhJ�
���\����?����%���s6@���
���h�һY��%��dL1OK�q��S!�YH��ǐ�MW{��V&O��ОsY������u��j&:�m���( 9�������z��&D�p_f7_��%�+F��m���@h_��G\.p�bm��q�C��\��k�D��V�i�O����,�*b��4u*����Qx|e{"�g�d�^�:N�-�	�rkfJN c�RB�g���b��6W=\������?�y��\����IQ�ov��լ(LKs=o(�s;f��PKG
�]|��Q�G�1�%���$�ŉe�F����Hm����E�[�F�CG�U�,�XA^�3r�#��H
֑��G����?��bc�վ+�Wr��iA�#7���m������Q�B&/��u�=(Ԕ:�D� �2���M1�'rA��O������e���S����<����W�9�9��I�}��˺^_��s��"}�y_�h���6פ����_�Tx��=�����������y'G���R��uJ��k�}I�7��Π�k8�ޡ<D�l%�+�LU�N#9ˇ�4CJ0u���[�\�~a��W�1%z�R����S+�<:(��H������(?�iFiq\�}k~�(��<Ŕ��F���^oф�<[��cJJD�0����2��+fV Ⱥk@vR�E�!��q+,��\�'��ŀ.JD��8+Q�Zr�a|9J9��H�O�U��/���	*�wW�o���LY�9ٵ����۷����/��7�)H��7�U��Ʌ �n�%�zt�*�t��\v�Li>�`�f�S�!tġ��P����U�Z�x,­6q���� s�WC�>
��D�rUR4��_��M�'������ł���H�ɣ�LPӎ��lI��vG4�q�zP�`�9��i���Q��s�|������\S���xlDd�p�chq���&�l���4��+뚶ԅ|/v����:%(B�^�5N^bH�]l�m�(
�	������Y�e����g=f�� ?��gP�IK*��a�)9�b���.�.�b@�'C���U��-�=��irգ����G����Ŀ?pׇ��" �2�ּ�An#\շN�iY��sS'�v؞����B�y'������ZI��E/	ț�\m���8�֛H�#]@���2��л%;�U�A����!�g������i�t��R-��M	�WV$�wcT��|�߰<�+O�`�a
�V��n�?�iq}H}[�V�yi���Ki�~�;�OfQ�N�#��_��Xr6�]�%���&��E� ���\#�X"Ϻ�(9�Y�w�YGa�d�� '�纚�u[�������D���͕lt)�3S�T�?=,��t5�@�=RM��9�2r���0z+T'˚Q��3�C�^8}ü:m�'}gP�%�kнe}r�� �������	x���1��?R�Xe>te�9���J���:	������;�~r�GC,I3O���J�/pe�p�p� '�A ��U�>I)��@h�/QW��s��O�mq����Ud9pS<��V�t\�06"��:���������UF{,�&�Go�l;��F}���5��$�/�r|4K�w��],�}Q�j�M�sG)N�����5���V�R��u��t���څqm���͹/
Su�*��Im�Y_J)�A�����O��2���h�_ea�ވ��Pt��4�+Y`��tk����X˘��l{JIoF#����MT��J`f���1���BW�1��������d!�]Xw�R�i��@7��Vq2ދ�oT O�OF����I]���5d��*���Oh�d��N�Q�*v0�=q�L'�V�\���S���~�;V^}a�2e:=|�&{'pd	#RN�Zٻ��p�p�(��
�=hY"�I�q2�2��z����5]����(�׫ґ���`�^��X��;#!�r 1;�e�Bw ���#) ��T��B�O��(�)3Z��xo7T�d�e�:(y��E�S���}�Y�\ӐC
w����J����n��X���#��D�1A�Dz,:�a�б���C�|Aي���ٽ��Cv��<84����f/َ�>��i���?����ړA:g��4�SV�U�<s����j;���"�M��uf��@a.k
I�z���X}� ����y���;���EY�d�{V��z�J�ޡʃ��sҏ/�>��� 1'g��"�p��)�%i\\�чnd�z`�Vn[��f�˵H��$.`��⽳�d���Lj��\���� �w��
I�C쐗,_1� `�s3W-?�d��'1�g���oH�c<�L�������.x�9Vh��U��i�l���R97>�?)g�,�^�3�?�D.����<y�/��� �;5�|Q���Q��<�Ao��+}nX�!�!��{l���s|��������\�[R��U�+>��ݣ�M3e 2�E�9�q#jJ�8�����`���?h�8��-[���<�tZN��D�sg�-@�ko�{���n8/�p8ִ3+C,�A�.&��C�[iHDW�&���	�N��[�ZL�"C��֫���{�&;f�W�l���	i�R޶�ڻ]�6<��SǨ�Y�L=ȯ?��=˃�U`hͫL�c�cX`�ρ��cJ�]��YPө����6�2��ԛɡal$V,�\˥�@٥\IvXW�����B	��� �P�2��A����"�.��*Պ���<��O��0	���{��.������Q9�������/
I*=S���.7�&���ݑBQB���֙"����)��.|��+?9�@"{@~)�L/���E쑅v���!ە��%��IR�k` �1��������؆�"���}r��͟���n%�h�˩@KM�o1�&�z�v�������.,L���k�N/�&%��F��4���H�P�*��.���#���\ԟc'���Jf>1���>��\�c�ޢ:�./�ؼ���L�\%��)�@�:K�~<:t���oP���~�t��fC��U���䚥7OG��:�dm���5.����ׇ& $!w*�w����hk�5�[$�[s�X�e��q�eT�'�J�>g��:�*z�������,s����j颗���f��S$��(D�w�f2H�-$R�;fZ/Ȑ��z^7���Ŷ(�tFܔ~J$Ʉ$�K�ІϺ��f��h�vש�
�|�q��C9Kx�ePY;�a �*���]&�P.��j|�`�ɬ����tтSJ8��s���;�jװ�Ơ�|+���Wk��ĸ��O�8���ͷ��L�ڒ��ύ�����`����g��'M�!���|;@�>s>�okmv��r�����K^�c+q�ݝ�Hl���1�	���\�h���$R����2=g�T����HGb/��6!Cf[�=h���Q���	}�U���1��M��#�}�F�Y��g(���\l���'� q};Xx�~)�h������>����s���90�=��Z?�Q���-x&����nU��Z��� ��I�n+KQp��`cE������c�h@���;��G�����<�B=(��V�����A�,i+�� }kH�/��t	��vu��ҽSt���y乜��u��D�]G�~#�ڙKl�%��[gh�<�z�f��x� y���Ab��d���CV`�����c����.���ti�2)��k�6���Ǻhj�#t�%�(��g�*fz��	�l.�9���Ϩ.�D�°�!Cؐ�Ճ-�����l~���^+"�e:�`I����6E�7(U��B�V���*�p>W���ݭZ����pw��*�@]JR3(�rߒo����ʬc�W�a)��;Y&�����h)�fޖى�t�fd�t���	#}�݊�$���)�M����0�J>,����ɗ1���+��54G�7�̇r'������+����J%�;��N��g��C3zQ�v�DerM�6�g�c���67\�(j�yΛ��d(h�u�A�s�� l8�wjji����˙9�v��l	�BM�?@���@��E"�U�M�a�J��A�ٳ�i�7�+�l��d:x���<�c!I�}��Ϸ���'@PT�����KUy�2���)���(�;� 	#B,J��俖�5F\*�;p.��"�C�k�N�� �3h�]�����x	��0գ�a��2XoDb;���RzM!*օ�Q���y�'|KwLb%h��ŝP#4�x����4���UN�.W�c��z.�: ��5h�R�8]#�5�?D�<~����X�@'���9)��Ӎ�P��6��MQQ'l���7�Ȉ�!�
����bHЩ��I�I�k�dt�|��,Z���C���/�W2i���$f�у'؇��_�P� E�#C���+��2g^DP�������3@ԩ<nK����z�DPf~eR�Z�4�
oI&�nX��˻��޼�qs��|&U�FdV��qcpM��*MnO���N@7�2-/F�^��q8�&m�S&*Ǽ�:sdO}W�`����!�Y��@�>Z��IO�e�x�gU ���h%b!�v�X�,��Z���>^��?�r0�0��6�gۜ�����e�@(D+ͷ�W����r�%�櫛[J�S��vc�����G�[��8��$�(�]�?1w�sSD���"`��7:����3��BW҅,)��$���¿�Ԡ200�MH�*�U�uWI�j���ٛ 8���p�0<�3��8o�#�QӾ&p��Y}���j�:�=B^Қ�j'�ڒ���f��4{�de�N��I�:(O[����`$�<`E!ѫ��#�	���,?.��/���~���h<XG�]�d�T�ۓQ��R��왎�Jݛ�=�9 �b��k\P.�y�Raņ�:1���a��#�G��[=Są8>)u3�l�grEJZ>����J��R��a�NVK��SA;�?�J\�urb�`z��_�9"�]޳�nRx5?�NR�� Ur�Z5�k%�>
rw���c\��#���/��Q@���٣���Ö����»���e�T���&h�pY�v,�N�����D'4��G%r,�!�׻�)sH<Bmh̎ ��H��#�%6X���_��2�O��\hp���~��+��Kө�'t���`���t�.Z����B�Q�Ʀ{�r��B)0O�8�}�%V����p+>=W�KvhəM�Ӭ�97��7*@m�i��]3�Y˹�w|Y��	dy�t�<�t�k�$��>B*��q��ni�1U���9^�
�߮H�V0�u�P��$;J^�pvħ;r&���Ъ	��w�q9�;�u?�˒8�V�
��\'�Ԯ�E�%��bX�ZA�V����ـSEo݁yœ�dNB�ȏ./�`C�*k ����e9T����@KW�M�����k�Ϊ�����9f�W;��*�"�Q��N(�&�>}��؎v����Ê���-L٩븭�c���^�qM`�{ ��-�Pd�����+�ge���{���7�X55���yE����'6���I�J Nb�"� ��zo��\��O�Ck����?.9�ZDr,��V6���|�K.Wd�2R.A9�p��>+>����HS�+G�l*j1P`�dNj��5ǋ*3�#�0��^(�|��"��}�=��[J������<����Y#.��M���"�3YL�Xl4ˬ�؜�g�Og��*D�+"=R
���p+�y<2�x�T��~����l2�*}��\��/D������j�4���a�1�*��d^�i�K+�~�U����G��5chA�>�
�ݳŧ�$�p����?��Tk�
I�6D���d\�N�?U�����t�G�\_�;�C�������E$���aN%�B}��t�o8�J�n�(��d�}n�؈u~ހ�&^������\��x��>>ǐ%i�+9JY1
��m	6^���j��{dS�P��-�V� vQ�'[��Y�uA���ΙPa���w���u�?����q��#$-���Ą��7wx�CV���+��F<2ڸ���j\:+�,Muy����pP��Α΁<�=:ģɱ8",�^<����_�_~~R3����C��-'@2d#�p�q]C������h����.к����w����a��d�(�1<����YL�G��Uɧ���P��NCsg��	~�Z����z�����u����)٧�3ܹl��t���I�J���
�ͦϒ\���V����U?��,^���Vm�U����"�M���HG�m,}�C���$�L\��Y��/%���a���7͡S��̾Q���霍�hd�D��p~sO��0A�����Ҿm���e9�G�.ێ��sćU�l��}�zsG��be�!Z���&մ'?|��_zݐ5cK��A߽������FLט���v֌��#3�a���A�X�X�
�c�Q�7ԑ䢵�Wa�9��5eg��K4WQor�i^�J-p<��N�G�.+E1
��h�ۿ� sp�z�CW�j�7�WM�3l�%�tb-���J��'�rvbe~��)��ӳ��� �뱲C�,��I����ը5�7 ���j()�弗߶%S8PZo�៚�᧞�V��ǘ)�:�=U����V^{z�.����lpԍ��p}ӊ1\��A��k���֒�G��v⒔��T���,��i3�jԓ6�&�r=L�� �C^�������j���-1�˔|�������1P�:fXDQ��IǑd�3��I,�
�h4*�*#к�&�!J{��,D�[�/��3��o���v/���[(6-��;���v~��wh��t�|�V)�^�ao8#��z��DF�Z��o�܄ӂ����Z]�U(V��B�!J���\��=noƨ��6��>���wd1��h�6�X_���_uy__K`�Ŋ�o�Y�4�Z&	a�76�(Ω�k��QM���;�}�3i|x��%S��&`�嘏��)�t�=�v�t[���Y���Ժ �ڐ�G�C�6�2����4h5�������C��o��F� R��G�t�>k+=�Ө�k���{m��5��q���!������6_�kA��t� #��o��R(ɰ�`N�븹@�+�����aY��!я񏦚�?�N�n��c�td��!M}k�^Г'U�����V����kS������`�T΍FC�Nyl�WXu�$�4m�vJ��=dn܌�w�x�����{��s�QR�:�<n0h����@3�N���N�����3���M��C��,��t�	Fg��ñC<�����yP���h�r�:x��y�F]�{��q����.m_R�g���K���r�Axjy�d$������z������쑕�l옪A_� �cꕮ� &z�����
�ϑ��p�d���m�L�d��6�I����?{ow��/�3%���L���w+$��W����!y�S����rk3�C�������Yv�~Pe��.���A��;8K9x���bA�@�f���
�}c,���VR���-x3�Ե5�Yz��3��oU��0�������CIÒU:���oB��J���"O�^��ͰO�[��+];\�	?����|�Y�)�L7����)S{��ܷ7@�_�2;�\�]����J��)z��{��r��E�p�`���yX�Oہ!s\���::��_��cD7��j��l՜_ꌜj�
*2G)���̶�*[,߸Zvz��3P�֨5`C��*ɡ���M�>~|X4�å���@�k#��1�.#v�w!X�#+�s�ϫ\�o؏obk�~~?��,$?�F�+��_�o��+�'�7s%�ɾ�(CG)�J�{1w��6 $$KD�"Yo�>-�"���Z�U�о
��K��
j�d��Hdoȟ���(7~%Z7=�&Ɇ�6����C���OǃN$�>LL�+v0KuW3kd�k�I�[P����W�CS#M���o�mO�A�NN eԫʣ��jK���09��a~��X���^ZJ�KcrI+�*V��JH��#Y&;kXg���f��HA�Q�a��Ce�,�F��7���N�s��H'�� P"F��q&����v_U���TG8q��?�b��T�d��:.�D�u�`�lR�y�-ũ_P��z��D����͛��p~V]��)���(	�8\k�ݦ����!pW��gc�Y)�=�!���<��
�����r���
ۣ8�O	��A�u���3����Co	�[yjLj��f�s�X/IpgFg���B�7���+>_Kt���H����8BS G\zcx��d�3��������|�e����b�nk�'Ka֐��ny2�R�L�y������19�NY��4;b���2m�voDq�lv�C�U���~�gy��lr`EY17�Ƣ���g3Γᮤ�D�惫��}�C�XX/�	prv���J�9א|��$��mS7��a�����԰o<������;�h�4���	M�&6	�U���+i.sH	�7�dc��h�T����@&*� ���'X̦pX87��[R���:�Mx�fr��*�1��w
���S�T��v��1s���S�-a� B�V�-Q� aao !ԧ �f�����z�s��.���HU�d����
��X�b��$�9 ���f�%����4�x��E�:���ه��݋���;�E��#�h�>�G�]�z�(f�e���H@��zw����מ�w��1��=�ӊ��;��=���"�I�b1�:vb����T������~(�YH}��l�X]��ڻ��׳\q��.j��V����W�*�I��lλ���F��މ��k���En����r��l,3��O����ϊD粘:�������@���"��"4c��Z���Ì���ȶ���γI |�bl��8r�cE�[\�Z�.�0���E�Ű�TN�����ڄ\�����7��ɤ��z�'؟��s��G+q[3�`�:u?Z"��P�5���V ����_���~�����kh9��l�j���*N󯵰�o(wҔ�m�p�u[؁����uv��5�)�dB7?b��bF�!�eJS�9��]!R;��ʁ����A9���ډn��g��l��3"!���􆤏؈�軶����V�-��������~�t�6��޲GΫ㼳�T-m���<��i+d�������]���d�r~���.|>\2%�pc��Zɶ�ڳbd�\6~'�U��}���nb������'�eT~�����@-Q�^{���oܸ7C.��d��{o��U���~���LZ��tq ��(�� �B�Ď�O�Y����E��N��l�������t`�%,��]+��Q�f8T�0x�f��`u�%��d�����V�	���`�q�Q�w%7�:��?6*���U���%^��DT��w��6�n��l!�&:ߌ���*�r��o��Q����q�<	1.W�:�R۵� �l���RJ��ѱ��߻�p�e�)��;ަ��GÄ"��0���P���vM�&��a���z�*3��3ڤ�编K"���$)����aY�b���	%�G�~�yA��fT@�}�n&%�9����m�6����E�F�wTV���Ƕ=�S?E��o�@�?̹c�%��iV��>��Fb�W\=���<֗ ׃@xp��[�� ���{#g�tꎡ���7<*��ߎ��
�v�5qR���N�h�M W�S�Ca�4�x��\^j���j�v\���+!�,d����\�s��,�T��J�
j7�Cm�vA���juw~���
֓�-=D� ���Ig 	��x�ȿW,�՗�'��Gi��:,�+@
q�����@3D˙�b\��p�� ?�c=��э�A	0c����%�C��@V3;;uTV3�2�ڊh��i��lj{�cǴ��K�P;��
�F`R�i|���������T)�b��b����ni�X��pƕ���N�xP&�A�����<��f)�L�_:��74� ��'�O��/?���� zM��B�3'��tvf�|'�u�� 8nIٵw��m=$�����Z��L[���Gh>5�sKP{2U��mQ+�F��~^j傱�����`'��yܩ�0�4-3v��ʽf<���O��e��7�d�qV�sQ(�j9`�[G�t��ƶ��W�����4�m�� �����%Ң��:'�U$����坎#-��Y�W�0�1Q��+x�xY�U�-<��D��e��4�,�/�}�YL㨽����k��c�[�S�%��͹׺k��Ds�4Ī��fx?�3E4�5�_W��Mp�XcC��֒E4�r���=e�n�XiT�nm�]��7�֘AG��5���VH���w" �#�c	�w������s4��|f �����1@��[Șc��ְC�vՍ�?�
�Ul���&���p7���k��8:�Kװ�g���(|���I�ǲ��lO�� �ڍ�������LbY��t�,�2:bi_��dgF���@�ystK�����X�r�r�L���`�~]8������!���T��Z\�>���`A���CnUk`�Dʾ��`o�D���S�['�а�jDB�C�B71����y�n�=	��Q����߿νJ'\�ð��C����Ա<�{��M?���X�9�7����K�����c��J�E�4�]t����o�bkս)_��t���4�9�E��|ɗ땪�ʎK"�
����ɲE��;���IRVL2=�"��?e�댣�X#K��� �m	��u~�_CԺ�"��W�`��pf�n�=|�:�q?LGS���EӖ*-͓V쫣���A�<�W�.�� N/)�v/O7��s.v�}�n08������	�r�`X�&R�6-�3*��߱V�5�Av@���he�Jy5���2�=b[���):?�x&��Ռ=��\٠�16\7���T�{u�4v�\eZ?��d�(2G�{�.m�y$s�_r6�ُ:�)U���vh��o�Xe/6�+d���+��d�aor��h��5V�u���~��'�`P�9� NTjo�,�E4�B̺Wx3N�K�q�zG)��cs-�"�|���cOɿ��ym�9�*.�E�m'�TR:6�P~t��Ed_��ER���{'ao�ڃr��%}ٚx0�'���LM�oP�3��I����VQ��h�l/C�[�R�����9���}Q+|�u�p��f��'��i$o�?J�?���fm���c���͒�?��(���t��@ spk&]��d�B#�i+)�ˊ%�|¼J���?YVyJs�AϚ;�&�9T Iș_�n�&�n�|�6�k[h���4�3�*#�������JWh�F�����Է�(!@�-7G1f��/�/GXO��GT.�ռ�Id)?B|��P���7׶J�m�)�ʞ�/�,�\�:j�i�B>GW�*ϓ&u��#09G��ioN� ��J!�����PGL����.K%�*�O+f_�"P�!Ï�7������������c�R���|�� �Y٨D�-�.3��

o�F*�&�Δ���`5+���g�K�U۶1��'!�?$��R�C���С�񼋓�*�$<�
H�JjD4�.xb�W�>)W��xtJ������OI�WF
22�.#�w�2��q�"-�lW�E�=�$�@���t�I[�ǥ9����1T9�=��>��W5�I�u  =���1�߼�(8��U�~6�^�ps��4�  x�"��(H�g�y��ە�9_ �ڛ~ŨnpZM�V
ʲ^n�Tio.��f��>��h�^�RG>�7>�[�{gΓMY��n��X!GJ�.)�D�J5뺻-�G�~��E��8���n�bV���F�eb%콚�t֡��k���ʿ��1ZE"��+}�����9TZN�UB5�F{��e9J!����8�C2���7�4}	ڜo\ZG)�����CZgp7����v��D��6�1�����Φ��Q�l���`�͛�g�V����q^�gw��M�2�� �H�<Э��x�m��/jD��s�:Nć��D�=0NG� ���t�3
�G�e�Ky#`�,ćݔ�޴�ĭ�^��ͨ��]��E_`�7��,���Z	�&��4��C؂�}N3��!�������%R�Cˈ*1�%ж��-х��{O��=�H�P��SŒ���6��v��wi�mbLd5K�
[94��;J��$���{�+�l�z,l:'crK��}-9��3�u+���-6Y���
�f���6�}3)3��{��ݎk�Y�S�j�{�|P:=(S�<N�9`MGq��X�~��]��q����R�ޮ:g�.���h�t�.�~��M��N�a�4���Ȩ����K��4����#"�>�^5�~Ғ1�g�~�������k�O��N[�����L #�q00d���\�>�,1f��:,}M��O�1?0������5����g�I��yH 0�)`��Z���,��t��9�S7�s��C������}�\/������Lo�$&s�N��ktkF�9�b�d���96��|g����Q�����ݲ(K��S���Ohs��o��`��,=�l�Q2g�񊯦�8�Qv^=������%� J!�ںH/�4�:e�;Qp�W9@�ɓC�[e��׫�+! V�D��� �Z��2�z3B	_�;	��7'��c?	CD4�g�o**οͬ���\h�e��g1���/������Qê>��l���[�b�N�f�6�C��V�%)f x>{ҿ=�5���KB�T)̩=�Ks�4~ۋ]�ñ��X�<�Ö��TU5�e2wu4��V�X�����2��3�f�����qf�-��g��P��@���F��dt�0�,7�f�\!j-�4��:�X!&m��ia��� }�HLJ��3E�f7J��w8��s#�U!����;N�s��"Zĵ�O2�m(�I������I�R9=�7�_a�dR8��!�8_�1��;r󚇷O-���P�n��ى=F��i��$���q���+9�fq���|4��1�$�\U��sQ��Tײ�0+,K�1eqrr�+A��Sk�����@��^	5Cnc��R��2���U��������E�$Nj.\~�L�U�����jM�"�� 4�K�9��Cer��^�we��bz���)ӮR�Vra���^���{o�Cfu|G94������Uꛢ��u�Z�����z�BU@ْ��峒쯑�W3�>Y�w��	�<��4B��:�=߂(�p�������[ĩ�@ ���`.z9�#�H�c�!v���Kx>Q0�^��>���&� ���c�ܾ|'_Z$UA�~	�����>+xԤRc����H��A��-�501����|^���R��"�t�G#
����A����(#w��~I�:x�#�bv��f�r������&�!���C��%K�9����x;@����sl�^�[kǿ[X��\[;�Avz�F�g�-P�ձ1򬢕�%�0���M�
>h���j��Q0����'/��� o�1c)*�i�gϟ��ݒ���P�������USlғ�1|�'v�=�륫�+�~Y�~�r8zn�ƹ�����,���
����]��Gxܫ#����1qO<)�{��J����B�E7/�X��#���0�Q�:)��]�+w|:@~�=��I
X�7E3�CA0�v�ٞ�W0��D��mʥ�i���`�(�u�V�X�G����3��j^��bp��{����|�:� q/��T����]��#��B/������6L^��c�*B��æi1�x��	7w�I�Hli*�#��i����a�-�Px����(<����\VC5��
�ē;�[vIRF�Bކ��S�,��lM��Ⱦ[H/�a�qXD����^݂�s�Nʳ�b����^s��%q�ԍ�$�)����xQ���R@&|�irmGm���X�O[�O7���D�{��c���׆_Wd�F�U�Z�����qȈ��d��v�vlr���)a����_%ɑ�����#�L�f.����x:x��T�P��d;����3Hޑ�W&~Z�%k���B tf�����l�1��R�2��\sa� "�LF�Ŋ����avw��(wDWx��E�H���v���W9,���̟��#�7E�yʢu���z��a�@
�)*��fl«{��iC1�8��D=���v����N�����+��S�� h���n�ƺ�k��k[9�r`0�8�>1��ӦSF4�|�-�^!E����+&� Sf�M�&����|lH��!ܪg��y�����|�V���.e<�O�	9�9��Q�<3cT�j�(��R�N6�:�ݑ�.��#$���|�����!�v�L]Y<�l|P�6�@I�D>�u�~}������)���/���M�du���A捵}����K� .�u3��V��鄯�����cP�w���*걢f{j�68uf���9�0A[�
зe�ysC���׉iv�s��$��� ���X���K3��.���)FﰝU��x��c�[?EI��UK�&���Ɋ���˱�������,w&x�cΦ�d|�Y	tt�5�D�HjȻ�c(���Y~��S}K�P�B�����_�'ot�{y
Mt�ܳ�m��!�9���2�#V�����c���T�3���ԯG�O��:��Tq˝߭ ��<;�����'p�}��\����+}濯
�I�/=!����n�LV^	o7�GK7��b�,�t�z�{N�sx~�p=�Z����7��?�k�Z�����/�2[�� 8�|L�Z���Z��7�i�xb�O�s���E�s$��Ȳ@�P��k��wJ�2�����Օ��Z���i������܂�$,��S�a��q�]�T=�(Z�i���F�C����I��n=�0�n! �$�+�+d�UO��eq��������ZJ8��@����n-�<�V,�;aÿw =�R�� -K����)yo;�q����R�
UF-H�(�.�M�vu�m���fh�g���*�`F�����
�����R�]ɫ���S���=|ĠrIܠ$�!O׵aC:��93I���j�P(mG�t�ƻi}h�4n���ڄ�z���e{��f�$:���)�e��3�Lriv^QK�'Kw����8�q��g���y�p��m�}����|��o����� ˇ2(��"��l��.%!7d��}"x� ���Vf�<����3��m��][Qծ9�Xc�JZ�(�*kv���Jm��no��&�������vs�D}�'X:,�z��9P��"���9W�a��p�g`!Q`��� X�y-C�aQ�k*��g�b����E�YQ���sNCwdj���,h��O|� ��'{m��L.ݏ
p�'Lq=�9��W`���rj鰕�J�*]%���[��Ώ�$Y%�ߖ�Vmu������� ���biV�>�\�l�NU��e�L8�y�Q�9�޾�&u%jyȯj�.���!���;�E�/&޴�Z�ޯ5�U�s���}0�cd� H^�~�L |rRo�j�No6S�Til�!CD�����b�c��D�䂿~M[��~�����3�E	��i-8�����?Ι���ſ2�c�������&�=��E��^^�_���s����j��UܥK����aK�j��Q�L��a��k�5��#c�ο��/�i�͹x�����"t8�oĥ�B�
��6���fOR�Ȳ���{�@-�7��t�Q:1�Y�+Ө��0���񾚵g{ʛ#H\�7�og���6���S����W"���wIjC�|��vC$�x�x��7���2cU|Y��^��)q�ym� ����ip�K/����u�������°�d��&+�f��AYou^��ɋ��F�+�"7O��ʌ�EZ0��J [:����z�f�-HMh���z�?���F�%�2�^�fY�_EX�#��#��{߷�	ܭ��@�x��/S%Q4���+j�UK�1eu8��D���ò�gγ���>�cR/y-�m���zÕ�(W�q�׿��=��Cf��)g��\��}���{�Q�}��IM�A�f��IQK�����imKYr��+<nq#��v��i��g� ۀрD���o�ӡm�ʐ3�ü)��71ܵ����:Ғ�rb�����%��M+	^p�\�""�C2(]}���"MF'䢬���N;�Is^q
�#�N]���{AyQ%�9�ٟ�>euN���%gW�豂����������HC�v�mU��R�4=�Rp^�Z�}��ȹ�	�b��J�Y���l�@����C�An�{'�'8&E�G��M]�p�L��BN�oԁ�B�T,UDt�R�Ǟ0>h�:I�5?A<��	��n�(��^�K�
JMʉZ�Ţ
j�f3����
2���n�v"K�x��s��R��ȯf���#>z�>s�Wrl8���	������}
�u��M���@g��]�./�X�eaݢ�ӣ��u�=��w��o���g&&鐯^�D���;qJ�'n�
3J	�o�̢ȡ����r��� �Г��J�DB��ƈ��L~ĲKJ��&��b}S �Y�°��{���t���X�\dٖ���3���A'�͗b�/6�랯7�3��E���\3{�����FP8��Yj_8�����?٦�e\͑ՠ@�gf�c��j'����[O�:�T�7�D���-�ćU'F����G�����Nά���)"����y�G�h�\�\&�����W7����=�*�aŜu��Ƅ�t;c趼��
��~��^T%���Qm��f%����P>W�Pð�mv�eO��*
��щ�pP;Q�?3�u��~�����,����ER"i�_�d���_��!��ธ}�-C�_��[��ؕ%���O���FFק�R+��n�9��Ӛ,+kP(��;�˱|Db�}��p��-3�[/�f..c
�b9��$�x��Ze*�)���f��y�E&w-��?���}/��VН�ܼߐ"�X�g#�H�9Vw��Ֆ?K3��yI���|���"k\Џ>���/J+��~�"3���2��z^v6k_P��c߬9�ù1��&�ǉ�H�7l�#��M>˰uihngo~Z�q��Rmť
�( =�-<�K���n*!���饛�!$���zRF�"�ۋ����7�-'i�N,�a=�Ir�ju���^؞�O3�e�_x- O�O�lC$O)F��)��`�e������Eֻ5c2���N�V7K+�Ã貤��Q�N6���h�F���٣&aFIT\�@��r���P�㔼�K.I�3�rE��� F�׊F���Jb?� � dvT@�6j� U�C����ٟcǖ�&2�2.8�X���&!�gj-O�"�o��J�j��< Ub�g�$�)6�Y� ��?��ьNN�z�jq�ָ��lC��b�K,T��?����S&:��^p��~	j��b۲�sIR
��ͼ�d,zA'���L����P/,�&���W����(!���}�<pZN�~�8zJ�Bvl�����B��ĳ)�����	��8� *�q���W9e�j�m���A�S��$���N��5 �.�����X�͙'�2Uq`��	aɲ�֪Z�"���9�|r�|�4�u���8�(������e�I8�;�Ŵt��-Lr:2��e�����>����$�Woh������V*П�9a�����& ��*�3��g���6���`���-��MJmOFp��ܬ�X ���r0�N��`��R��;q����&����Nī~B9Y<��F��^9T�2fso��g*�@*3A�j�SI�{.�wϷ���
� qiWC	���xx\�p=!	I"�p�)�'����_8�a���EE�
�.�L��BHHS��n�HY����:)^����Zv�����j[a&��z9�<J�.�c`q}���u�X+Ǎ�OLEl�.v'n��A~�?��0]�f��}��'�j ����n\<�*+�Z�y�*��G��(q3@.C�[�?S<�ݷb�6�m6�/,�b�q��F1��gǻ�m�s�Uo�G����_.� .&�;mꯛ�s��N�t�T?,z��#�f����5g��l�L�����'e�ꜸѢ�7ն��Ü���(29��ּ^���$����F�ȃ���(]���K�|.������b��2M��Ѷ{��:4�>���f�*$Y�!\	t;jY�(KلK6s��y�1͹��Ri=E��X�o�������pb��A���Hr)X����5T�&ܨ���'�u�L!H���!��R㷍H�d����������ͱ.�H?������Y���~�Okœ���2x,A
���ع8��uB���gk1�׮r��6�R��%m<aϏ&}��s|�?3g�E0����8=��Zڏ8X�鞫%���qW���|�A{�Uh���ψ�v^�6P�N]s�I8Q��q�& �
c)44e��'�^*8�D�< b7��� �G�wvʋ%�E�+;͟G�@=w��tDϘ k�,��T;��'k�.��.���$�,�=V�]��"�w���C>�R�i0ؖ�����öz=�/Lp_�a�fHΧ�e'��鈷Я\D//bR:y��*{Yg���V,�[��w�=�A$�9�,I�p~��q���`�ʣ7�p]��~j�ߍ�P�#Q�� �e��E��i�tϬݺw \�xט�5s�x\LZ(�ѯ�s�$� ��?L����O��Ze��0�����5<ؑ�i��fK��n���2t5RN���~㺍��Ql�� ����;��[�����p��L ��r�~+�����B='�����P���� ��F|ݱ����z>�[7C�׹����0��ȍɓB!�n�o�2��Ed���4�*��ʵ�ɥW�tu  O
q���ȋ6I�Z��}H�7:�宐�����{�_d2��>\���b���U��P�-Z��|L��0M2Z���[�,D& ����SV�@k���r����&���(Q�FB�ivp,�c
���/���sM��͎��E�B%g�-3�	���GR�XX8��~�NG��pVy�y�$r��U|9w�H4!''��V0Nj�"�H~p}�d&i����9�(Ea�4�yy�k��qr��-�<P""����@�Z針�P:RS �tx��2�����gN����(Rzb@0_
� g�fJ��A���W������c�����ڹ�����FG���]?A�&�]��=]z���$_-��3aY!�F�4�H�)��^��FeRnэ��	�+/ѓ�C������;�x���ki{�_�m9vv���1*]q�w�*�aD4p��"��A������MJ(i��B?)�?����1�����-���ӝd��MG/�V��N�\�ũUX�KR>��*����N��7{�	uy��:�U|��~���s���&�1\Pt:��k��f-�I$:`-yw�%�2j3�C�,G�;�5���qU������0����N�Q���Ӑ��UzNl~E&֢h��]�Z>����gB�[]��C	��+�6�4wYͿ?M��R���k�4�9v�c�7%�7M����3)R|����D*h�Vp�r�&�hiɶ�3<��|�*lZc�D�,������}�y��`�R�  �pjK��-
�b�,�vV`�à���WUU=�֡'W5	���Qָ������M@p��n�ĵ'V���_tqQ�(<5�}�x7Ul��kӡ��i�X��u_�+��o��~ɞ���dZ1�2����9�5,1I׼te�S��$4`�O����\��V� 	q�3?("�mҩ�o>��ΙhӺ>rOZR��`0�����qV�.��H]aK�l}��s?l�S�$MWq:�P���]"k��L{W��C�<�$�ݎ��B�x}����%�O���h�b����Ϟ���v��>tVuw��x\Y%�t�au�����[)-��}�2�y\= ��y]�6n;YN�>$��盙1,�?`���������`��	f$ա�ϗ^���Ika��'����΋P��gi���@,�1!����� �%A�
}���OB��{���_��0���ga0�7u�./UE;���Թ��~�s�
��W'+���)��)#l-���:��*��V��?
�nrm��B�zJo����.�+}b(͠���(s8m#�ѓ�T��C�h���>�PA�d[X�_u��}�Zv�خ���{�*8f�缐���>7�\Z穐�5aʹ�W��R#�r�4u��z�J��&҂�M���n��ę>�� ��Fǿ��֥VJj�v�!S��+
�œcs���B�`oX���%Dz�,�AhK&�S�w��8����{����7cQ@�_�W����!ْ�T7?�p��m2uH�Mу�gjf&�, �#��Glm?�� \������h�Ƙ��W�Ȫk����������{8������(p�^�
�D.f �3#���sTJ�:Z+�N}�#�s7�JB!s�����]V��ND`�2B��`b�ƧZ�~��z�P��Ltd_y���'�����19S 0�?Гp���!�n���̅���V�tw�".�1�6��A�'^�.�ڂ��BpZ����@LM�<���i��6::��~�kFo��:k�!�����$;�}h�=�(*���4!�W��cA���
�|�� "[Q6 �S	 �,Y���sf}Ŵ�0�!V�7v�9';�V�v���b��Y5q8�f,g��aԏ-qÎ��'9���L׫����皱Nzs{<�bDJǻ�q�����J�z��Y�U|cZ,���s��Bt_�B o�TP�J{m1�L`'8]��o��U�y8m���}�'�Z��L�"��8�\�t���5j1=��]��ʬc����A�^�����z{&z8��x����gZM3����'��i�T�׋�w�nc�;����9�`e`x%�2�ȑ����0/{dC�7#���w&�dJ���,�G����i���87��tuR�N]��� 0ۈ��]��d	5���4���/Ћ��<��x��ڥ��c&\ʉ�Yu<c�f�Rl����������J�	� �;{mx�1�O\Ϲ{�;w�ں���J���~�c�|��;�G�[�+W�����X.��$��^Z�4�U�l�\TuSq�3sSj���O����5ֿ�)�D�~��F�֚��P��uA����86�~�XP�	��Ҡ$[V�!g��3U���ͅ����)3�	����nzV8�T�#;�V�ߵ��e�*l�sߦ��l�t6�Gpp��OHr�L���(Һ,�E�8 ���^�[Oݤ�[fC7ĖP�r��4�.4Z��5��3�#��j�,�*ĭi]�9�l�ߞ:m���E�e�CN�����|Չ%��=����B��^>������GIb�=��:*;&��˺4��\'ވ�?�Ӫ�փ�7��+\�kC'���.��Q���P��B�_�
��F���ږIߙ�b��I�m��>X剟D�&�z`4�۟���H�=Tv�[�H�����d��Û����y	�UNڎ:q�=�h�G�0ۿ��K��6�\gi6ێ����<9��98Qb9%�5Z��O? P��(��t��4�]�(:�,��׍"�YY����T�J>��m!h'jz�a:�e(�U>���ڄ��fhosi���Wuqxɤ`���λK�Zv���Ǯƶ9v�Ί�Rn����/n�\Z�D�?���*�Y�.���T��U�ذ%"�Ό.��t,Ln!���
w̔/�&S1v:דJ)�+�~�:d��m�Ǻ����m������������N󨙄��TZ�cz0��J���;"��Gg���|d\i5fI͓�( �h��B�J����0���V�JP�`���!�����
n�n6�ş�џ�@���^�YQ4�3�,�����W`V.$91P��W��1L<*�
�/�yox��V֮�����@.�W��Iٛ�1IؤoI�Gݭ�����D��[����iBO�R�E(MW����Q3��4�h�=1V�'�hg	P�Z�/~�Y%ШrE��sl�2�p�ٮ���@�?�u��X��>�2vj��	ȝ�i=�}��vH��= �@��]cb�/a��r��-A�Ҿ�ﻳ!5@�T��si�!j����"����������ë��F���o�8@`���۟��R¹��k�,G���HA�!�[����P&��AP����Ǔ�K�R��u���3�uD�=�#S�F
�������%k�����<3?�>��V��A�Iw@�Ά�Ȥ0�g����v��Ww���灿D;&�GOWe��9WR� g��h��!���R�A��D�NhҰ��6߻�uTW�z`q"�oC��º�<�����E`D����x=�73sRC�h���6|�=�e����jI���m�e�ݩ�ᔩY�>JU{/{˱m��$; >�/yy'u���F�/a�A=�cʸ}�m��6%x\A�������~�r;>NC̃:��!p����X۞��+wp�FF�����Wǵ�q����Ԥ.�3c����'I�Wh����I�ny�x��E:��{O�-��歰ӷ�̠Iş��X	�K���WV�k�r7:z�V����������G(�g��v�j+�T]�}��	F~FP�X�ձ���z���1-�m�@n�:q_�P�.�U�z\{>��#h�ڢ)F
 ,c�1��u2������#���C�o���]����ᝂܛ]I�4�G �`�%#�?�g�Z	�ئ����hYi��Y%�0�g����8[�!������PŜc��'_�X�d"��ӫ�\a�8�̜�r��1�s���鳝[�5��
Ȧ50;�@I*�@�c��aqHlu�b"	�T�"e�5u��I�oV9K�B���R˕�N��������	 ���0ᅈb���C��X��`}�LrK�x1��~ H��jz��P�q�Ѽ�q�r8i�a�PB�nV��@7��V<�Fa��t��Y��V�#�:e/�_�(w2����\�e���׫ǃl	8;<#ྛ-!#����D��1" ˊ)�*��W���!��5Sb��_z��s�� ��8��m��Q%(h�;�<����O�fǞ�~v=��z��9�:=Ff�m�-�������+�x�!��(Ĕ���x�M�tvCE�}�{3�:���=�07`�^�(Ni�+Z=G�)9�>lQ����ۈ���wIa����m�I��,���
᠅W��L~�&��ogL�l?AR����W��8�D^���[/��L�Y��
b�d ;$G� %�|B���^����$�K*�:s�(I:fUB,��<9��;V,�P_]3s,_\�*͊ӒF��^אt]:ڼ yA��
�%չ,�;إ[�xҞ
����
Oh�t�ܢ�mzwC�&"|���<����"�f2��Mp����j����z�-��A���,2d��{Q5���+��t�kX�Ʈ���1~h�#ȵE�H��Z�y7.Q}
�g���Yk�m��K�\�_��OZ�I.�;�R��d�b�lj[3I��#���Ð���6�9�����L��wֳ,A���޷�簑����!B���%g\~CK���E��Ǔ����&���l���	��+�r��/���Z�cm�?ނ[�˖�L-`"�aGc�*G[rY�������;��֍�4yK�����;���/M�Z�q�z�� 0��2D"���<"�=��Q���˅,�bK˩Fl�^5 ?�<��/$��{�A�C����X��"�XI�Ϩ��ɮ4 �Io/�O��}CtR;��TF�o�����%��	�w�@2j��&�!�d�=}ur������l�b@g�4�����&����=xR~Ϥޅ8y�D>�{×�'���W��bd:�.��7X����8CБ�8�}�\}z�s�+U=<�
��8x��QY��ꤽ���x�ʠ��&ST$�y�Rf]��D�~Z}�^�@�QN8y���s<}Kq��y� �>/Od{>7H��li�D=mꛏ�i�0Z�S�8�Y�S~�*�5"��B����iU�w���5{Y��3��U�x��ŋ��a���e�� ;��j�o\%�<���,�%�۪vp���K�Wr��a�@1-۶/QP]� %{n���M�m@��S���*̭>e,�So�{E/�Α���9.c��wEVӋϓ��{W=�#<_���� �Y����Ա��ט?�gK���w��<n��e��3�Gⷌ,�NO~�zz�����sDI����{���Jw�@~M7��Aô*��S�@@��j5RH�|���+,�&�=�t_��p�/����]#c�-JQdYG8���G�-��OD��AZ�*մu�l�CN�K�zm��+�] N*���㏓Aцo)Q�{-zճ�"\
���'i�9E�p-��)�M�nQ��bb�Y�����o��V�cdq�2�(�ʍ�H��pwkz��)�EĦ�.Ř{�PD'	.�!����А�l�;N�� �H2�8�����ܴ����V��M�r. �\j��3��e'�(��Gu�у���S��Č?>vė�p�͵����$���Y�z��q�7d��`�S�1m�R�Q��_|��MA�'ou���j��ROR�����`.E�"u�/�X��*`G�U8&+D@�t���!.+?��c��w
y7�jO�H���n�ΰ��EV [��T>D����N��r r���p7XC}���kc�mQJ����x�5]� \^���y�|u@�G������:*;���3*e���o�;����m��3��(xQ��1�H�!8O��|�t�F�v�Ă�V����fz@_�a��~G}�o}�����o�dK�ح��ٙq���c�K��`eø�\��&�~ū?;>�D�e�j�!�zb��[�Vx�vLB��-o��`��	�3����W%w�/�z���(i|�A�
�r
|/�c���קy(YY��	˱LɓH+v!�n�|;������'\�k�����CZĘ ]�(����)&.��^�;��c�����)�����x�xϤ��B����> D�4}�S��`/��dݒ����n�[>� ���=�w���#��ZP�x>N*2��nR�d�	�cH*�.kR�OP����oҎ�
M2��Y緐pd�7��ݐ	���0�O�Bޘ���@���F���Eg�dW�V��F�����'��S �xVQ��ϐl����";��T��R�~�1k���n�I�t�	/�/��} �/��]�I*"���2I�J��1��U/���wRK��?��:Cm�R�W���V��J���.J����ϖ���_^��mt�����:��1��:���LO�Cұ�I#7�m��z�8֨7���9�,�8�!N��֦ܨOA��<]R��dxh>}l����v�g�C���1�KAü, ձ:C��S�^�C�#R4������h��zcN"��&v'��
��l�"�DhWؾ�<T`���Ã�f�9!���ǚ��W����U{h������#�_~��'j#�t��
�y���7��+\�[���ڜ�R�2]�'��]ޡ�S���݄�������)z�#�g� $�r��OSǧ�v���ր-�D��m	5(T���B*8D�C� z��^�ڦ�Kz&�
�?��3��d�¹詫�=X�EJDA�-���n�T+J�;)���?�;��y��H-����Sj���+�b��^�BP����@ӗ��<h���|��H��,%�(������{(�WP��{������������E�z�����uM��+�x�T cSH.?<+����O.	z4�RS�ǐ�G�U�1$�l*QQ-�fs}W �m�Nᢟ>������	��������(ɓV�»��q��ҼXJ�����~�������.��LZLC�@ف�K|�赕o:w\�M��O0�,9�+h:C���5>,�Jb�Rv��Q�	��a�$xؖ �}�y�@�k�R�ODb�"�2Ǘ��0('��{	�Y�|`��9�>V�r��C�������)9�;�����N�<�l���<ԋ�$<QnۖRp�Sw3�*}k����5��/�he��n�[槢�q�oP�9I~Ar�趾֜�=�qL��.�T��4)���j�c�?���}Z(���0&b���%�ֲ+PPsJR\G�9�VP�vv�mOs��f7�*o�Z����+���V�b�����K��Nm�-y�}7Pi�,�?��\h2�0�
��C���������l�J�֋'�����)@\�F�A��|ԛ���R��݉c��T��f��ص��H��4�d��&�o� <lY�]����L�)�]{D��)�N� D|IQd�0)�9Ї��=�ű3\r��T�X������B����ΈReɩ��V3[�g#����C	��ǻ6X� � �wv�6} �����Tݶ%#7H���������]53���\�Z�p�?Ѿl�F�@��Z��
�9W��p+>!�9h^Lc�x�����@9Ku�_9r��ݺ����RM+�M��?}�!Ԭ���������s��7�Ա��ʚ!��.�R������W�^�%��K+���9`{f+��1+Α���Gk���ڂi@�4^�V2NX�� SR�Z��S�!<}��X��nG�_F��3p��f�����қ�*���tNCe�5��6�w�@�d�����q�D-L�$.D�� ˖0� ���x��^����&�sb��}h"�Q��-zG!��e42���yF���{Bv+��d����icmA���SZ�'���n��Z0Čy�Q&���7wp	g� ^��[�+����Z�i�D��n�"���9���!٥�I�_N���-���z���(!�/T�?�A.����;Kȸ&ӥKG"��4!USH���f��h������}(ƻM����;K����KY���XP��	j�Z}{��H�A�Z����m*φ�
ġ��hp���h�:�<[n�w�z~f��Z͖���G=wpTEc���<R
5�++�7���R6�T�M��'���g��xdͶ��]Ć�����y����4$[	d�yh(��WQ�qmr\���A�r\��ڹ:)��t�)+�ܭJW���I^H�D߼-�\.�璉�j�ш��9�V4L �sz���`7��Ǟ"�*0sX�=-$J&V�.C��0e�Vp���A�Ա�'��h��}*�$_l��YӲ����g��S>x��-M�T��fW��hj�z�X`Y݂����B�+�kmn�5�9�M���9;l�je2�2\*�Y���I�-̱��M�h}S�|T�Lph��
�[V�݂9�n�d%�X{3 ��[Ď��ߨl(P(��A�SX�x�t���� ��R������F�|K��K��''�]A傝9������Oůa%{*��
N�=K+���6Y?[��"a���{�.
ALt�Dh���q�k!A�|����J�(����^-o��x� �N��f���z�����Af��Y�V��������<���ԯ� �����ϰSR�ůr���cJ'�� C80�� ޲��� ǾF+�[�v'��zz�(`�Hۆ���_�ͪ�#GmH��ՔuI����@Ui�U�c��v/���w��2UY�
�Af���2��
�2Ks�2�4�K�"��"�
Rʍ�p�5I�I�:��>��N��+�nD���m�n�L*�~i�+��@&�4YY���]9�� ���G��
m�fc�DDJ�*1i���N�"9��4z�i�Ňg��⋛.�}��u�J��b}X�Gܟ��ϲ0�³1l9��zF:0��k�}ƤGVD��k�`\K�k3��0�.�/�N-ћ}F�$��&���n����b�^�H�[vF��a�ˆ��;����h:.<R�,5���r��_E��TN�?����Xҙoj�Də��B�#�	�'���<�A
���D[M��i_a�.&�z� T�[-���f�B�R-�Mf1ɤPS�iQ���n��w��P�rR�����ؠ����a�b�x������eXy���'�ڛk�@�4�N���S���d���~ȳ����A��^�i�~�J�B���$��% �	�$�\�e�wHG��N��d�9�����8S�I>A�ѹ�4C�%3���o�ױbc���)��)&�[��u�樍v�I�aoS!M4y�Y�i�Jb59�М�br5oJo���ލ�(7At<���$T�{�F�����9�&���ʴ�e9�='t�ŵ��U����t@�U���Fn&��4ǔ0̣S�k��-p�}a�L��X�ݛq��dc��'nB��q�u�8�أU����z1^O��#��R�ϋtKڇ��i��2ǨU ;E
N!۰ݲ]%��IՅy`��MS�*Pz=nɧ������o_lSX1��Cc�*\�<������\�g���}�t�T�:7��a�[��t���|F�L�"Gn�����R���+�.��PNۗwW�w"������Ō�\��.�H�ŀX7ݪ"���ɱ�{5&J
��uɪݍ)�f�,��>����1�D�-h�FB�ț�Ͳfa��p�M*�ۀ\sT4�S��O绌�L�h��*��J}5���=J�8='�*�n=����ӤEx�Q�衮"Q�A`����Ȗ��5�Yo��~\��
��\R�cpz�)�~���Q�Ѱ�mݵ8�B1�h{׸"��]^��[r�����'��_ �`(�C�3	�'�Q��f*��ӑ���n{1��n��0<;'B�4�qȴ��M����Q��=8�/�)V؛����� �Vg��u��HA�~�E�Q�@���n�*il5��{H�ZV"��,C��s�/����`�Q�kL�5C��(�Ω=�h)^}�iFr���Ԡgc�Jz�:rs1��6�� 4쇑(yB�0i.���P�V3���Sd�es��=��%3�rq���عC �_�����X�E�v�o��/���!ɱ�~�)}�߭X�.��>�5잝�I<��g�(��M���J��
��/�����V��߲�[��s&Z>�
�� +J����wc�+t_~��"SO���S�=]~S[��"�i�L(�e�]�Ֆ�5�T���菾W�N'���J��CJ�~�GU-���X�G#k��x���	Пɵ#r�m冔2Iq��jƎ��f<o`�g�h���,״oia��Ov�Ѻ�&��hQ�_�������R��&v���}�W��i#~��X�j�Sq�s��>�N�6�M��5���b;8z���#��E��%����Ѓ��.�X���.M��:���'��	�:�u�y�{�q��t��E��G��j;;�,�����bTJ�����L$��G���:��L3��l+��b_%��8j�V��o�z�9g�������.pc��Q��2���V��d!+��(� Z �\��y*@�Z�Ee�f���s�Zp,�ݽ�3�,	��2�{}���Ü�-�3>�%X���3ue�cQӫ>`�a��G���$�;?-�X�j5!t�i��\l�Y���H�TCUڪm��ߵ	��i�x����K���W��̚1qcF�{���`[2�^�g\��IH�d6�~͒T"�"��L8�г4w�����W%h]gdP�]�X�M|�iH���ofo' �mCE۩��sO��_1�6�n�:dڻ8��{�n	��O���{�������5��8;d�D�-���h6����h��v��Ӱ�;���jk�$�..b��&sR�8�����dPd���(a="�yn� �}���H��$���>�A�ǦU>'���v�,_�G�Za 9ZU�8� h�*�{��5�FP|ӣWq_�Os_��ܖ�����f�K��nZ[E�� ���`�����Pr���O{�U�����ˋ��˾{�6	���@F��`���tX��d���tG�2,�t��o���%Jm�6<�o��f��%Է,�=�٤��R/�Z�n��w�z1�NT�mv��7fp.�|VU(u�T��dm_d{�JY{�TX�
�}�T����}�>*b�y��J�L�{Xa��#G��I��:x��	>��`2�mb��V�՟��ܱ)~����� uA`-�7�na����Ӕ���mx]��������O���,�	��dGxÃ�b��YWqIz	�����usa_�]I4�Di$�'~�]���K�����x�.�ي�A��"Ln�7�-|B�:-��!R���Ou���G��)�.	°G��}�B���-���ޝ�!���;4Q������l6сO�I����.�*�-��
���|�]U��%8��P���]���܊u&x�8X{�F�آ�%CM����/s^w����7��`iЛ<?�d�ɼ�x=�M�d�kv�5 y�$��	�S�H�(�x�|τ?�<܀R\�}��7��gM���]pr���I�r]��ML�)AcAAv��P�_�zf_�,!�UO:2Æ;���G�MOּ���y�hƔӀ�/=�E�W���L�T#`��u���#���L�7����H<ٰ1'��P���	d���j}���䀳�_Z�w�nO��쪽�`A�7�I3[�n�:�>��Sg���/Z\r���ܳ]�2�x	R���b%R���h�u��:]r�^��=an�G$���!D���
���n����崆��Yd.����*q�b��(ʝecm%m2Q1��ά�VcL�D�gL�2����M��SC��kNX�R�V�̼ցgUz���1�{�׌t�fdwU����j��ޣ�4�\�\IL5�x�r
NPϖ	�`[��!�	���|��o�v$�4:�FB�*/����[P��O���p�8�C���na˟�����b��u���i�PRo��.Þ�f��b}��i��a9�e�)�7��=�&�ejDcufG-}�@��ÒV��l�a�G���䧴.\�d�Χ�������/��+,
���]�i�ʃ�$3x��5��^Vÿ�+dų��wx��9�\68
�;0{� ੎� ��PH,8��$G�}��B�/����~u����ݛ�$$�+�a+?��T!b�D;ݍI�듑�^����f�C���Z�� ��
3h-���	1n��c��r�s�<p,dP*���9���u�ݒ_/G�K��'�@r'�&����
_fh��<o5�J�o��*ħo���T̸ޠ�hզA��
�{VE���0߽5��0r�F()(�����!����g�P���;FS�󖂸DK���-0�47��{Aj ��?�Ij�3S�Z.q����h��$�����\�D���}1'g��ld����-�oA�]�g��!6C�؏*h�+x��W��n��G�b�mv&%�K�� %�:W�f�R��at%5��iĬE�m^u�O�������^��͌��k,���&ێL��E��Dϲ[�H��ޑX񅳄|��s��ۇ���*�%EزH�S�"%b���V�f�a?Mw��cS���� ���)9��?�VUl�G�!=];)rFR0�7��à/$���	�U"���B�N*a��!��#�*L���8�����KZp@�~C�|"��w����S�7��̝e6qi>2k0�.�A��LNU	t�Y�w����՝�`DT���*,�6��޵6Z,"^U	���`�nmi7�A ��G���DW����� i=� gY/Q�X���l���sF�8�З���f�̆9�b��ԥ�?�R����߻�z�;��:&�	�ӑ�Ra�NP̟'����H�:nQ�CtL�n��⟣Qa�*!p���%٤n��L>����k�n4��^t�~�t%ydj]E�n$ V���1_�]#��C#o�7�ޢ -��u�G��ǘ���ژ:���M�ʒ�`�pj����p~�:��X�&��
Y�u@T�+�/@�wD�X��^�X�˽l�O�򫳹�]9�a;Ld�Ԛ��Nf��dF��K_�>� ��A������K�],x]X����?����$R�Ds�^y[�^1}9AG�V���ti�tu����.$�2�����AMdL���}�FZʖ]i�U��+!J�7�Z-�~U��	�:�9���Ɣ����P�E�d*���l�J�h�t�r~+.��y���2يF���Z1��`$�"@f���]�[�	�;vx�0��̩h�m�(�Z_0��l����U?n�ѐs]
�Ϯ�1��M6k��J!yV�e~��f7�cY��A%��RP�f�s�5K�h��]����X�1՝s���gD�P�56�//�`�0@���߳�[9�_���^,��?Ϛ�fBB��_%�Mz�B}�$�Zs�ǰf���=�遛/H�|汓al��qo�]�l��b@H�'\��Gzg��ilۈBk�R �EN"8j����)U�3�g^�t���>L��E�O����7g�W�Yz�'�G�fd{]�
Cz���t�^*	�
���d�!��^�~�����Α�b]85�Q#���)�,8$��p<��]�3	1 ��=��`UmƇ�r�z��g���t��s�;���t9�f^�㚻i	mS���Mr��jϷT�[J)��������uu
���7.Z�Gy��>�9�tI*���(!�>i��C 3B��=��a�����؋��r
�V�0 jY����8�u�Ø:�:�B��e�~�EP�c��R�j�]˥9�*t�m������B�����8��n|�Hm���(� 5�"��B���O����p�ZD�r�=�/8)�D�Q��q���6c�,�^m;7�;���p�-��/Ҽ� �P'�p�T��F9��X~)�աc^
�D㚟o#���!��������G^D�&�G���G]':�ň��agP�sv�y��W���f6x�����W�Ν�f�z�����ER�L䍥��Y�?D�8���%}�£���S�V���P�e�9����rTe���f��%�㽫�q}��AUhҙ�뛳�֖���F�H����������b���rQ��E����P��A�qǆ]��/���7�
x:ПRl�x�7��d��P�K*�5�����_�0��8-������Zp�\��f&S�Y���}�o�@��ƱŌ�y)��'_���/�&N
��dck�nZ��=�Umt�;�{A"���M��e�r�'uVS�PFs����2��OE��l�1��_ѐ`��]a�#�������`%!�J$��
%)N��I���el��U}��)h�s,T�(�kci�Z�2����ք�o�r��)� '��(�'���=�;�)�B\��!���Df<�/�W�T#��7�UL䎮��W�J5|����g4�����������ب��s��t��jo\v�#�w@Td(Nib��De��?xX%����L#�;����ܮШ����:�e&����J<�1uuR�!�μX���"�!�b�����lLy����}׫(��^�>f�.6�O���-�?a|�k՟�%�U  6�Z�ؿJGN�������m�(�`�GMY�?��d\��D�\!�M �Ϭ�i�M@Q�`�Q��vP���Wg��r���$�x$���o1E8�v��$W��৔`�5��"�sm�R
�����씘1�_�/���~��M�T��Uz����3_� �$�=�Xݔ��.�$��Z�pJ���������`'Xy�<�b0҆@��9���]G�;�o��`�A�3�>JI�Z�"��#�y�'H�)�p�D��?]��e���&�T4�'��&�c�#�#��wH��0g������{ևz���z�3<��+a��RvS�����O�1�zĭ���X�E}]f������d�+cc�E ��,h���N:-:�L��D4�"��)	)���c�5�>&�T�`kX`u���w9 C�/�Q�i�����-a&�2D��`#-��.
:�ܐ5ׯ���htǼ��3٨�!�p՛w��"���R�^���n�Ӽ?�r��L�T|L�BՀI�i�ڱv,�;��t5�	��$Ag�����S�ȁ^i������6H��+-P���N�5��V�SD;l5� Ӣ���gYһ����؛B���ׂ��<��%yw�7x���Af
ep��o��$���R�J�]-2�u�n ���qk4|a�]�����l0�"��i0�D�s�e|�"�Y:l���vF�	ѽ�x��q��"��_1YՒ�qn��-���@yB��"��MU�ނ��0�R<��{�~I�ꁋ�s��z���M�a���_��0t)�;�q�$QW��7�e;W�����vƟU�E�-�Y���SG��5Ä�j�pD{u��[>�<<�_7cEDy��X����q�f�{d��o���6*���&�	tz���}�0��t���P�y�%6��4w���9�F0����D_��ϡ�j���/�v��gqH�ӝ�@��`j��3�nc��/�g٪�ζi`zl6�
)1{N�Y�o=e�8;�ˊ�%إ]ј��#��L�wH�ayk��2fu��O�L�\�Ͽ\�x(�!�['��e�V/R-��l���F��>OL�;�~�+?�l��ɍ�a�	�ī3Q���V�s��]���4 `R��ØͥSn��)�˕9�&�+����HdF���2�]���b�<��7��������l�<>�m�'�JY%���tL�G��r��~�
�q
1x���
��T9l�;�_�c���)u�ǰq��g� Z6��+�u��`�E��,���w�e���v���ݘ +[�:J�d�ry&|��Ҽ����L��]K\��#�7�*Fl!iJ@kɺs�~r{���E��U�Tf<�����P]��M��.0���<c%��Ք�]�.G!L���q�����(>�6��?�4]��2|�w��F_5%'��v�`I��Ô-Q��>�+Y�����>�k�?kN�u��Y5r#q������
jݠC����^�y����*p�����	75�l:��o+��Q�Ad��+�� 4�Kǀ64f0��Ȓ��|C�R
�[J�	Ӷ0�gud99+�~���
��[��}'�?���R�a��(��3������2���%P��M��N�'���H��D�gB)&R��*���%Ʀ�J�~�A�{V����L���	�ykO��B�g��ce�C\��^�9���︄G��iW�p���K��3ı#��
�S��P��/1v�H{�es�Q�4y�v	Ի�[V��#�R����<���쨜6��B�&~��Κ���F�iR��5s5�� T� "�#��!| C�2���j9ϟbr8��&P��/U�dy5�;hᠰm����sJm�z�	��͞���*.�̜�02�º�vi�2H"�(��T��=4��ƚ�n�� +m!#�����E�isoAjA�t��"DY�PJހ�o��9#+������
e�D;�3���������]j��i�"��n����ty��UД��)追�����aB�D(�s�a 96�΢�<t���ksu�����YA�=*'|����δ�R����(,�,�Qfؽ�<�C��\�������:�[5��<��/֔U���^�#x����������s�5]� jW��E�G�\���N�A�(�Ao�SCQk��|��֒Gݐ�e%^HV��1�=l�}���%6�)\�e�ayp�N~3N��1��l�r��p��$;��B�SȺ/HRZ��.իf�Wl�GX�پ�ڎ,����eX�D[�|����)_�4�W����Z8����}������ΠY��/�L�Q�sc騐4��ض�	��?=_��n�����3����w'��g�_2���z��L����q����K�\�l_ƝR�勩"��7C#�0�+AvH,�jy[�˫�Lm}����$�6^���`�q�5͸f�����
e��j�:���HM�5��S��r��b�yS��|.���w��H��pK8,s*g�i��Ǘ�����7�5�msanƥ}Ï��<#�e�(>^᤹Qgs�X��@?a�B�S��K�����m�f�>%�!O�D��E�u�a�ⲹ�h�Z�� �L��{$��4�fб�=��#6� S�Q�z�ϥV�*P��.c�
d2Gi���d(Һ��sq��Ji���i}�����ek�J3�U�Zw�b�i�>���c��v�d���-<>�D�o*_�?�-�᝞��ar��Sݫ<eG�m,=��z<[`�R��=ɯ�5_\Ӷ��ؾ�6�	�[*8��Q_�>�7ʞ�Q?y7�;�ad���ן��Ux���1�1$� ƾ 8{��{��͉�dNat����3�j�����A������7�%}���HW��e�?�� %`�{E����LY�]k�-HX�����Ӟ�ɭ8B��^�+���s��_>���|u�T��$�X�#:^�zɜ��5}�a��&���]b��栙���\��`��W{E�DE��Wճ��8�AuIu~�K���mQ!�/Q����S�m���Y������,�Z��c�jK�j.ƕ?}�u�*���������۽I��a<�d�n	�-\�(�6!�+��"����Z�٭��=�����=&�VȥXB"��%2@��f؆�I�qr@k�B�ٛ��;���z�%����K�qpe3�0�K����Z}4C��#�Z
�#V��A�|&� �?1��tȸ�k�M28Xǿ��5�V?���1�{8B�q�N�H�k�D��b��݋<\�2潒�Зk#��bB��"�G�D�5�C���w[SX} N�7L#?�۰�#a�p�s�X撿Z .����}�P	9H�q{�C�"�?pEiz\"�.��H���&#����1=��f�|�gc��9�갿V�9L�|+�΋����	�_������xs*2K�Cī;k�-�CkQZ=�)T�(����0�Z���D��ƻ����:��Plj�Qb7z�[�;�vՂ�L�����_��ܑ!�&�OmC*=W�#$�T�<(�-�Ł����
�1*
�tըA�4��	���:�sc��j_���n]<�
�%p]"a���|��EI���X{j��9S. `�>.{�C*������1F��^�L8g��0	 ��6�VFAO�AE� �3Q�������H�E��g�������L�M�/Ep$"�FV�> 4�h@���q~��ZNY�%6̭�כ/�i�����!����'Ig��U6�aÂ��dkN1v�ܾ�c���H��vc�'���v�XH�L��v�Q1��~ҥ��|����&�R�!���H4,@42: �$�}����t�P�O�\�&�w���2���C6�ɰ(4T{*y�{0������{�)%x���8��{
O�����
9݀�\�Q{�GRT�3�a�5x0�!G�P��o���$�,���G�V��L��ϐ�r,�I��Wp�Kş�>�c��N`سh)�/�$�[ζoJr�(=@PΊh��>n �����R�F�B��_R�;Dd�r/�%����5��I�壋�~G>BK�5����² [�G�5�}��R���O={JKr���[�/�)t���j��}�5�Ԑ����a��*sio�Z�%9�B�CF�m��}4Ž� �$B�M��5j�[��M�ea��L������T�֎
"K19�ӾA���x���5g���w6d)@]��_�ൈpG��ʝ�1�ۓ��~��*m ������wgM�<�@��P �[�"���cK�� �	C�Z�r&�wЉ�+b�p3�[r m/0Ę/�QO���â�}����֦�8`�3�y�9����}�*>�9]$�$r@���8oj�?f���s��~�|�KU9�ۍ���r�R��o�Y�WFN�tG�:��k��h߇;�7�h	Xv"f�֭1ץR��ڭ����t	��K���Ξ�����#)���;b�.U	�>4��S�xx]�sU��q[����k���0ߘ��R���.[�<�BFL�������;�wm�T�k�i�s��J�"CB�)H�;�FTr�[-GUՋ0�@H��z��#���#��rY��}p$�R&ER�	$zn������x-��~� ��f�4eCl���V3
�|�0�ٹ�C�(�A�:"�l���!�p�
8�L͞��e�h���pD{��F�u�J� �X&j�!78�gn����N�]����C#���2"CW:��9|T�o�|�/�6�z�BX��%���0�Ji�;�P��+�_+�i�/�v�!����m����	¾�;+9	FQ%���}kIe�>��'�TV��DX���μ
j]-r:��۲4�yEL��4��'�� q�HFBkӋϚk����I�P�q(J����)�]s�j���"d�����@^;�;2����P9����x
a��y��{�C�h��ṥc[Р��>�zP|����R[W*��/./�����h�g0���[��ݹ1ٿ��8H����bAq�NUnK�%�,�g����Ptc�:O
q��["|"�`��\�:��tuG����#�/Q�rKS}�JW���f��w�L�X�B�+��	?n���,����Xf�Y?�xϸ��>��5Y�lw�U��R�R>�1)C&�3���ce\e�m�wb�1&�=@;3|r ��R��4�@{�O�=~~���3{l/6�5��� 7�1��[@>c�dל����;����*hS��#���z����:��$^z�_�|�)rqp�"��]�	�.�����%#�9M`�b/;�T��%��|���R�S9������_����#x���	_���^{��h���kHߍoAz7��Z��H��:[1`W>$u��y�����X���S>��; N£�D���'�[���GВ�O�b������X|D����n���W����� PX��l��$�"(���rb�Ʈ�.��C#��'�[��kї�����p���)��b�&xRg�� [����г�ʖ���FY�Y��;{�g>���f�c?�`w��Iw����Nu�in��+m��\����a�y�I�Rf^�'3���?j+�a_$�6E��Eɤ|&k���V�~���#���0�|�$$|�k��΂	ͣ��ݔ�J�2
���ipBi���9�!�(�dh;��(F��.V��T�9�!��Kя.Y�{�����ҟ�8gY�M���t�ћ�ݲ������"��r�]�9��qT_��k?�K���0Q��/Z���X�n����b�V�uD��e���g�'N�H_'N �Z�G�|��0�@>����]$��p����1���Rg\��.þ9�"!�*��BqU<B���1��Z�	��t�Ln��^?jV��T�;X����l]��46��d�����,Y��kv����XW����ҝU��ҷ�S���n7c'_;�2�O%�3�����'��ۺbH�]QR$C"��z�
�1)��4�J>���@��N�Zeh�1�c���X}��]�ߢ� N7Q'��F@��[�4+ ��$xF-���(<�A��c���F�x-�g��B��¹�7��Q��*J� Xt�������+�����(��E�s4�	@�!��Չ���KJ�W���6����cei"�
X��-r}�/�7'�YH���0���ß�r�\�N,2���UQ�.UOf�ze��/ �W�U6# q�1���[�샣���� ����_z�Ȗz`?���P ��t>��3&|�3�t�V�Za�&��1����'�������N��/Ln�[A
�B�)� &]���Z�o����0�w��#��M��/
�	O����ćP������)*]G��RMj��E�G��{'�N7��.1$R뀕�NƔY�~�����[�n�8w��q!?�Wq��gT3�fB{a	�ʁ�S-ZL�B����/���Z��^l�]��}�S�j6~޻q��ڌMT-�u�r��(������H��K�D�������.K�t%uc�H?��Z �����qκTt���T����0�<V�L��:�[(Y�+@t.�_{��_��>+f_�����'�x;Cx�|!�*����t{�wb¬m������0�^)w@�Ӷ��0��#|�d��xĀ�:�X�v�[�XYa���V�gZSjb�����4_�w\��G�Z*�DI��k�/�Jp&���s·`��$�:Ke1�W�c�ςi=R�ڂ��d��Q�;'	���J�?j".	 p1�|L
�nv��j)��K'�Dc�m� :���7�\���Ge�[��6"<�온3�-�$)O�sz�w ��9�"�m�u���g��Z�q4#�t��~�"�m����P����,߫����iV��E8�W���͊./�b���f��������Ci�l)��M/mXm�ݕ�{Y>K��E��0����&�(�I�M:�M�����|�+�5�a<.�P	���;�ſ��*�m<�_ȓ�CXf:�Y+��6�ʣ�De�֣���ZN��_K���;O���M��A��w �ɹE~������ۮ����;����6F5C�J5���7ή"a���nݻpN����8���ޅ�h��x��6�����6��۝#m�y��3�VXV�������D$���6�T��m�%jJ����.��g��v#OxE^���`��K8�LI�͝�b���k�:����7��,�y��޹̑��q��f�z��n�_S�[̵�u��w��[�y��,������^0b윾��
L��L�zP��Ջ܂ֈ��C}���
��&(5��e�mB[�t�7���	L�S��9����ˠ�y1��gd�v�f5h���\��`��x��[�G-�"���)	�f�R	ͺ`�YI*�,�]�r]/a��oz@\��	W��Τ�?�a�/��'G�X�_�C>�ġ�u�u*6uzу(�TC{�xU!�'��M�[Y/�՝l:-����;�����ſ�K�oЪ6y��aDk�k�ﾹ��S]��5���K[�I;�)꠫�:�3)dzr�n}C߰�����f�#���û����P���9��=���ɨę
�6�q=��P��S��j�Yƣ@6-�U��ͼ<�#�#���$�����R������"�H���wʘ�.N���$V�SR{��7��Wm��g�S�Ja��H=!�4Dt�`�;@,��UP2D��
\��2(��豙�L�=���T8�C��6�2T�D�^�4���Q�Kn��8��L;�B�d8s��k�� ��~�6n�V�N9�y=vq#����O�Շ���aE+�\ۇ3�>���/�5Qz�#O���T�=~Gq�o�z]�P��K��Jő������<`ܞ��]�m���v	j�ڗ����C� ��鹭��i:���^���|�CL6�
E��?NԽ�D|�ן����������[��(��M&�蟲�8��0sC���uءH=�s���V|��O�]���$�6[ Zh�撀�]B�g^'�%�p ��O��W�"ƛ7�������o/�3���i].HM�j*��<v���v��p�uO���;��/m��sth�iC1�gM���:lVxYA�E�*�@�~��
�?�&�i�tŃ�K��p�zȹ��ۡG�G��lj;>&���pІ|�Y�8��;��N�+�$��q1?�"�;�NT�J� �~*<Oz���U����r�ړ�VU?c���{�\��I��hI�M��������ɓ#�w������
,h��cV��֦dd�F����;��#)�V�Yf�ZՅ�U�FrЦS��<mZ-��6��ɕ�U�����bmo�9>?�~�6��Z1���(��h;�V2�`.
�F�>U�<�q����]}#x6��BښiEeu��X�J�<b�J��x��
5��sPQj�V�������;&!�a����,���H5��۞��S�� �J�oCvȬ� Tޯ^�7�t/�����]&�D�L@0A�]�0�=T�q-W0�.#����eϋ�y�a'3�/0�̺�ϴ�Rv�D�M�:��븮���W�uD?<T�2�"�N�:�,����T�5��L E{��e%�Qb�~���bM�U���OR�|�,W��fҎ ^��2�
�#'��G�݉����I��∘�8Ǽ��=�I%͘R��w�4)�����K�Η��A��1g���Mm�rgV�vs�=6,�@�Ĳ�BU�>��_W��%�I�OÜ�)(\�u�΋���꼟X����;�-�������Hj�i8���wֽ���p\/�B�Ș��C|���S�8x7;{`m{-.��%g��&?�H�ɛq�M�T`��RϪ��"�+�Q� ��Rf|���M� `zkS(V��=�d޽��xD}0����&4��˨���lʩYZ��}���QNW״�
1�vs6)��1���.�JD��Q���=�8���0l��P�̎�'D��c~
1�����b��*�r&��O��}pqO��������'���+k��ތ���8������,b��e9@㯕:�R(��@�m�>��j�a��c%��j���!sn�^I +���o'LwJ=��ٮ�q��"��Z���]B�}��u=a����?�ѤMM둑-�?���A�X���L��L�~�d�p�(�v�f��ڑB�q8��6������.�� �q�y̬����F�ލ%؝.<4��F�P\Zw��~�y���5���4���
�U&�� ���i[��`��6d�i ��l�J�42��ɽ������.�ߪk�Y$�] <���Ie/��{�?����5>W��bq�#��4�q^�(��ӱ�����u�=��r1�SGp_H�Y�"�R������ur�msm�$G����;��:M�"�;U�.ք=.:)��������8���V�N9[�IϏ}��A�йaI�IΈG!J�c�{;�ni?�I{zF��OŶ2)���#�0u�x�i�k/	��A�t�q|��R����ߩm�S��a�?~��A1G��b�Ϭz���������O�@�,<��/�?Ԛ�� ����n@˭��6P<%�6t�2�Q��+����Pլ�2�/�h���g�ݕ��I]5��L/�y��Ŗv5{���D9��4������cJ�<m��-���5.�_v�A�����xK����W����͔�I5���Ps�<��)ͤ��Q{M��|�I����9Tc�:GU�j�E"\�y�
d�l��n붏���ч}��CQ��?����)1E?�j��9��U���蚐f�p4��
�J�aō�D�>%/i���ߗm�yi�7T�����8cA��/�1g,A�>��5y�t����.�dod��D��U)ؕ7]PJs�wV�x4;-�;�QӬ��J��o��E�d�O�@|�R�w� �W��j���/�V�v��DH
����[�Ď#y��PS�� �nx�n#ׅۤ���R-GJ������X��_��������lU�E�����QYt��~�4�Ĝ�U]�X��}u�[F������:{�/��~��^Ww���:��dY�B���B�͎���ڞ��][�١V*��i6��t'3�o��>2 ��B��^�������Č/�CR��bْp�t�!�1@��bU���z�t�sRJ~���f6LQ8�MhnGD��B{u�U���' �fO䂒 �?w+	@\836���^D�^��"����s��m�C�?``]�z��;�����_�'f���/L��S���Ƥ_�3����>��*� �rNQ¬@łpG$~���5��9���'��742�����d9�j�F�)��?�K�����Lwe`�B�����}��"ׅ_F�|�&/��� &�å�.���[��uv� 񳺽��a3��߳8�+��qX����e
h� XV]��w���n�K˙��K!�޴�{
U6Xܨlr<s״� 4��,�jr�r�؄�|�mgc������ậֽw@���X����J�n�G	�>H=�i�m2K:�����R� b�At.���Vk{�<gG�7���X�zF�}���	v����w&X\T4���ȷ";C��������/�.b��\�(�ԁr!��r���$[�cban࡙��jX��M\�}&k&$�I��=�%wۿr�u�V�α�0��l�����z�`�偐��/m���{"
d�_AC�ŋ�J�CgN�;�5���Ϩзy��q���	����ϿG���i��~�d(�{�O#&-��'t�� *�Sf�R���UM��3��@i"�P�/� �:�j��܀ɕ��wS:�g� ��B��"�p���X!j���0� Ȫ�Ѱ��?ْ������.�F�k�N_ ��)�����G�^�r�z&S�!�W�t`pV�SX�mF|��ȟ�i�,"<�1��`�/����,}"-~�c������qG��8�!�L^~�Ҕ�E�U:�pV�ZX���Z\ �" r�id��۶W��0<�.�_o>�W���.|���W�}��8[�7�3�y����i����n�Ԭ1z����`t$���8�ىT�}Z}�'�q�l,M��}���_ "G���g�\a^Я�J֢�'%�b��O��˼췑��)P��hX)��i��!�Qf�g&�v���w�8����,h{��W-�I�n�|� >0��c���g�&�)6����݄��h��lD�!9w����ۗ��O���������ͤpJeb�2�H�A�F�GQӼ�x��F��g?���N}T{�:^���?�#�SUP�:��N��\`��~�_E@��P��i�������E %C�֣i~�������+( ~&uSvf=�2&��Jx���@|��̫��`���"�I
!ߕ|���d�^r0�{�Oe|*�����>7"�ڒ�f�������{�S5���j �җ�6�A�w%�R�鵉hYd~��������)�/�$^�劶���_BpG�F��o�!�<�ϋR���\�mR����J��0̤��w����� ��+����9��]�wX`��[[�5��G/i�F8�.���������n:�j�(�vs@�  6n4��	�x;_�u��e#"�ZdB)v�S�솇J����'�(�|��G}h��Ԣ��9}<@���6:;v�����C��	�+|m�*�u�-^��a�������|���hI�J�v"����YŲכ��E@ݮt�\��d��փ[V8��p�i͑����2K�Q�%�@�<p �-@�-ϡ��^4U<�h
{�Jz���L��A{;Ψym�;�nV
#GT�&�MY�$�!�ڕ�3�o�'�q��l��V>�Gc�k�Q�k�����ae3�K�X��jsv0J�$0��è�(�oN��'^���Ю׹C+<�*S��#
ɉ؂���v>���n��^�$�2�׾1�U<|�2]Yw��{V�_r�BY$��^�ߍ����ϴD.�_�/R.�B�Ww�����j~o�/1R�iW�
���f�;�(�0\���!�*��Q�z�4�Y�h$AN٤"�T�l�lH.���O|>���h�CM�5S8����ꈢ�jsp��?��nV˰c˽%�s$���I�?8[�,g~��d�P+"F��>J����M�8t��")�8���@]��?1�4;���P�+���}��QX��zR].��lM�`tEȼ'�M����)`\}x_����lCCIA ��Fڜ���9@p��/���S��:{�էr�!n�y�3�\��ČJ���/^�z��3�	46���1"]�*LMmK���2�Ӵ��a&%R!=:<t�ƕ��!���6�z�m�w�	X�������EmB1a)$I#�(���l�f{;5��Ə��f���F��'����a�B���P ��k?�B��]�<��
  [�o+�9N�����+����̜8�!`#�6A"�g��x̼����6;��Ҷ������q��M��q��A�Ը6�$�c��]I����<�XV}���
F!#�+ۑg���;ۿ@��'t@q��q���)����h/�Zn,� F�^��C�}A��2n�+�M�-������ت�3!�C�׋_��7�yP�!N'���G�ּÝ���j�����é֍��ZF*j��ُˆ_����r�O� �Gj���z� ��t��ծ5ʶ�ݼ8���s?� H�Vf�pԫ���/%���V���[ۖb3�o-�&El/	����%�KJ*���̐�! 7��n�͡Fn4�c�W�zx�p7������?�uM����Dx���M��W�L	 +dO�$����Չ��i�cD��a����7�m�_�Y�-h��l����� �,�}�Ѕ.8�}G��ҟ&-�������@�'*�M��=���<SZ)�%a�?Q��������ڧA���t�!����>T��/,wm��P.�eS�3�L��az|�ȫ�r� �:;E��so���05�]-IQ?�%_M4��0xuU�Ԝi��U��W=z�`�$�Jc�K��VC�����(��֍#���Y���q���T�_Y/��z��X�n|�[�{fJ��h,�F9 ��F7~�!3@�*��~�KE��F⍜�U�}d��Dw£49Dm��\�� �+\y!���m�z�"��2��s�Uz�h���D�G�Jǩ
�_���:{33Z9~�Y�,TF��Օ�e�E�h0���� r�2����K;�{��Y�Zi�V����F� "�`�򧙏(AM�b	�"pz+| ��pJCf!\�C���"�W��@&�I�բ����{�ɻ6�>���R���b^�qat�QY���n&X�X�ˢM�ߗ���f����� �uQ��&l�n �2	�9*�a����f��6���d�]+J�[;μ�QE���6�B�*в�g&S���gXq��)Է)OP-Lt��P* x��3l���..���+�� �1�D���Vs�Q���L�#�?�m6n����8n�����)WY\����=6dE��$��������c|�iS�ߓ�7�D�����{�e�p�N��~q8���,��R�~�X���h�`�Hw+��h�:i�%��J�-N@-��l^����X �F���6��e���7\טB3�w�{�W� ���pJ��٥������{i�k�n..G�a7x��)�T���<�]{&A{��8�E#�eT�u�RL��������HW��@���K�9:N$�n��n���{U�����$�"��Eq^RM�*�Ru�WX�sr�V"-Z�ج�S��4�D�4p���\�U�yr���1�`�Q�n�q��E�+1��h�K_��;u�>�)�_u��F�F�r�w����g%s���	�Ssx���oFV�OL����H\�U�^��;�#�tu	���k�R���K��ű[�I�'�"��u|\�2yH����l�sC����'A���{��w���v���!<���fIx�0�t�
���JSۘ�p��^Mv7�����%���T/����Нt��?UL��;��|,/�c=�1L3����`�P��:4WZ]��挛 a��ʛEUea�Y�=� >=ۨ,���ؾ�VDMם����]��ȶ��%�Պ��?�J�GL.��8s@��%	ψ�ڐ��L����F�X�o_��X�Rb@�#�E��Ϧ�����Lޱ�\E�(�)���0cA���Zb���sb[Y�#:����:���8�g�;x�������i^�̓V�̊��AD�Ì�L��,�_PV-<��� � ��)����)�H��?z���.�ك_�1�3�\Q�	ۉ6��9��=�	�0Wy�$ͬ+ۃ����ܰ��q*+��)�v��/A>{/S�v��>�Z�[�|�$hm-��u9�$��&�@Q�/�� ���Z#��q5���4�VC�b`f3β�1�����7S�fQ�<u���BK{���E��(kTZ6H2�/������ؒ^G�������r�@E�4in'�g(�n���|�j�wIv<O
�O�I����d�9��My<#LY�E��u��D�R�F���z�p����0I��(���$�龞3�lOԇ��.��>��1������ߏf ���<K�|�&SӐ�� >P��1���ا�,e�6I�M��]lэ�Z,��/�����`:=(�;qؒT��,W;�Ԗ��/p����|���� Ѫ��S�
<6m2
�Q"�?*G���-9��c
��}��(�����9���±~,���F�͠�*�4�>Po�Iw�FN�E4ݼ;<;���[�k4aI�����%c9�ƽ	��%�����8�=y�Z�m�v#��$��]g4̽ܶ�� �S�d�}��g�wI�n٠�sׇ�\�H�<�T�0X�A(��q��QE�`�k|�6G��������|��wT����QF�L��Gg����U�����p9�9cU�F�Æ��
WђH����2ʮtV��힦����I�*��LWn3�Lt|<;ĩ�`��!~��b���J�
zN��-|ji�J��`�߮��G��^����&����C��_�m��=��!{�ͼSQϠ���P"���yo���?�����Ң���1�Cp��I�����٦�8��mY�W���,�c%ꜳh��J�u�Mb�4�5��N\�!��E��� Z.""]�*7�� |`g��u�%�^o���tO{Ek�)�6,��8����ar����m,L.�L{�s;9ۭ��b5�a0E�%4�������
0��x[�Ɓ�� v���4�U����� j<d���>��ě��p侟�n�*=!�_ݣ������b�-���ѵ}`YY�a��E�W��hzw���[�e���%Ƚ[a=>M��*���YJ��F�J�H^O����^|�Jsx�ͬ�/�?,Л%|&[mW�Eu�M~Es�o�u���.�����nkj�����}��"뗠n`��W���X����ʫ"�o�Rx��

Kol'|t.�b[�A�x�
n�b�_����s�:�^����Px�]w��ҝp�w9�C�ܹD���K��	�>��&�FA�Z��Ӏ�7��e���wr6D�ԙ ���\m/�H9�7��#�dѸ������v.ۙ`�<�=���oL�X8�UC�DR?��Ӣk�2{~\ͼ0�-�BR�7�s-<�4����Eb˯A5Y��C�8&��ы;sh�4��@#���`�D��%D#�@�(~���h>����m4��}��^`	����� Ȑ���csB�>�����Y�G&Z�tdE���Gi����Қ���������p�k�Z����JW�g`
�K%����n�����\~���Nn��#ky�_��oհ8{�mƶeS��)#�Hۘ���'Rh&�:��3�ەf�<�`��l�Uz@G��?�ef�b�E�L!���I�,�	�k-L3���UJd�]xVl6���b-�^�7�$�p8�"���Krkx�$��ە(���`#쭧�'[��I��)�Lk�y%�hJ��<�Wv6�������0�+�ι| �9�m�ɥ_��G8�^Nx����&K{��3�Ro4�ֵ\G@���2�k��g�"����"w�!KIj���J�[|H�S��D�:��9�P�.q�÷$���	� :����v��rFچmvp��ㆨ���S�fE�[�A��W7y�c�B�q�}5-?b����r�ؼa�AjvL����\fK�[�/g�s��
�tŶ��h��ͷ��_�˦`��
�d8��Q�a��+����0L�3���C�3�n��n��\Ƈ �fU�t�ӫμE˃Pս�r,F~�I���|��հv	]��ѹ����-���A�]���bQY���z	&�C8o��L:�c����^X�1��c��`oZ��A$9#�2�ihL�_�À��k���ΰ�Zh�g��Z�E��a,�������雎δ�WS�|-Vo�m,�)�4��j���[��b^~0��M��N?�{�]�B�^|KF��3���@�|��L���D[��JF�V9�Ǽ*��5Ԓ��B�U��͘.s�B�f?�͝�,x�[E����q4�5��f����F՟ȴ��fHZKvW�.�8JF�������+(�n~_G��4��Qi�f�C��9p�W{�M5r��MȀ���rnVz�RN덌r��k`�/b�����׫�8h�'y��w���RU�wv������Z,d-X��
{,	Isx�Y�-=��]��=�/Z�D]���Zo^��ƹA��&pt�^*ii��Y3�B!�͘�-��&�qZ*B����o�C���X�\2�t�Pp\ 5S7�_��j�ϸ����H>B\�t@L�a�wZ�"��bo7��_ܓ|Zen
�Ɣ��WГLkWZ������k�{�'��ꥈ31V�y�ȰsP	�g1RFg�VR�0��Xd����K�BOR�,��V3]~q�x�M�A��6W��t%�ʤY�h�`����Y1��B�kc�I��Gdi�v�xsh���߅6YB\):� h3���r >u`<d�Y��PA.-���{��$��\��|u�ؙ��#.S��"�ӟ�w��.DF�=gN�vم�\82~����e�y䝝�[�+�I���o��3R�����Q������\�� :��B� 垜����>�\VF����p0HVse�.k�b%�R{h%�w-/��v�1EX�α�,��(�1�G�X�"���>���~X�X�n^2M�i"���H�I��?A���FN �H	�c��`P+�` uo"<�1��6��.�|א���r��خj�?M%�_���̖S�7B�3�{���� Uc�m�~��
Y���٘�f��.I���>3t�wS�{�8�j�W�>��9EKn,'d�&p���Q��|��»܉l��Q�r�7A(��I�j� �6u��Ş�9��Ag��bk���ެ|�k<�qq�`�F�3-��%���=X������z��cD\�AU�3�B���m_CZ�eս��.w�y�&r�Ɔ2ߺdº�sb>v�S4�n��G4WN<�4�M��,$_�ەX�La�n���@Z�Z�3[�B�H��g���9՟%9IX�)���C�0�3P�?��
��!��ػ��R�:9em�r>/1�P�\&��
)G?�1�~�ǷZ}o�����6���6o�"�H��5rx�7�_���e��8���8�~��oU ���KY��k,-|H�=�0��6�ŷ��/ċ�l� �/� 8(9.ٟ(*���ָ����| �D�[n���]�����R쯲9�H�4����=:�(�<���2�����]��tdȠ>@��2A5�Ib;��' ���e��V�s\�*�� ���1�!����X�.b�ăn3�+�����YVؑ7V�|4���nE����Lz��x��bƤ���-�W��>�[���>�d������yi\�KO��0�Ga��E��[?�3�VE�~��a��H�w�"i|��� �c#�s���L��CTyTS�5@��7Y�"/Tn��<�+��W����q����h�N��ж�`G�����k�-�-��\n��w�:)�\���o�\�u:�a��#g��mI�i<z�~��'��КKu���S!����d�����Ia>�c��Q]!����10���S�sS���Jj��Jn�{��/�rd&��E�� \=��a�]�`q6�=�UM4o.�њ�W�0j�-l�
�<��~=�L�	�iP�^#�g�d��ƀ�D�����J���C?�p����k�D(|;�3X�<}Bg?�S[=8���i��=� ew�{�[�� ��Ru��\h<>C�E��m���х�D�i�+L�	����v��Y�)=�NcϺl�S8�̻�"�#:�V�����M�����FF���Ii ����h̊���Z>N}�l�����4�÷��g�y9C�O!}pk�b�j��h*΅$G%{g�z�7�U�GA�P}���H�Ȗi�
h�/��Cbd䝮��� �F杆���K���6�`m�F����|i�\Q���%d��晟���v����Y/�Nٓ���]�p݁󏑩>#SuIrg*���PB}��%xm�R6,���Ch�|�O�-ć�*���W��W���R"��c�X�5�V�Q���,�A}��2�s�	�ޘ�)7A�U�$�n3���/�.�J�Xl6��
a�f�u��D��҂��^wnQ��'5R�U�;W�>�/A,���l����B�>��U�i)t��y2
f�6�6x����X�f?baD��G%7Ԕ�T�5��*�2�=%?8��t`��N��,@��V�o
��t�V�6U�&t��H�ǁ��ȞQ��x��H�2�u�q�w�<�Wt���
x*ؒ�~�iՁ#)�h���Xm�/��?M�:L�!>lss3Q���8T"N�P� �C��> ʗ�5c���")�n���,���ʜ�Ͻ;q,�"��>du�H�#r6�:=�F8��>b$^��)Yb��˂j����z�eva.���|�����$�*�RD�8�sN�M�e�7�lX<���2�|�ό�9c��H0���f�Z��쉞�B��"8�a$	�z-�f�a��,�5V�uC�R��M�x���!鮼��A��箘{�u�r�L�/�Fu�4&O�<9��څR��]�(�L1�/6S�D��}��ѵKD/<٠��m��8�R��<	6N&|�K�Ua�c����ń�PDceN��o__aU�{v� �r�x#Iiy� M��p��[��:�$p G*�(��2���^aBFm��+z�B�iE����`�=�bH�Ӯp`I|�.�� �X�J���e?vL�CZ��5�{�E9?�LJuQ5�y4���� �}���x�z��l��E�Ig���s�d�d�1�r N��{�:������0\2�#�<��P����id����*V`^3�4�c�C
�NY�L!4m{�������Y�P��H6�1��})_�zV��uӠ�ʢ�´����F�g������;E��
Ø� %
Dg��k/��"B�0�7��v�G�U�}R�]�`�AiU���K��kA8�[ I&�o*)�h��J���nT�02��ąγA�>�uɄ�̒���.sG���*�_��e�UNP[89��$,��a=0/�>���j��_�$��p��Vq.�D*��.KG�ؕ��~�E�ɳ��8H�|�Q�ɛ�$�pܡ�x���4]{����Y��h|�<6I���]�i�����i��<�� 	9ZUk�� Z�GezԢ���,�Hu֗t������2:d7n'j��=�s�
.���c[V#[��BBfS��7W�	扑%�>�e�0��,�m>�H��\G����k>�+�^�c��������~е����XR"8�:+��80 � =jQT+�������M	���^��0��7��KB���k6฼c�'t�Bu䦯\6���X�j5���,�SS��x�`E�#Z��j�v�W'
8z	����CR*D}�0�j��{��i/_���n�I"�i�x^1�8W;� ����R�kd�� ����o �ǂV�u����Fl�m����r���p��ݧh	ǡ���O8n/YKzGQY�x���*���7��,�`�"M(
�W�q��L�I7�����s�R���(Β�P�Y9�^������4&w�u�ВoF<�y~�$�Ja����;�]d��&��!&�'U.�c��"6�sJ��Dm�i����e׏���<�]��v��Z�L��һ7r�I��&Ӱ�S#)5X��)��|� ��Zg�/[� ��=J��ZW������>,�����1�г�N]ߚP}*��ʖ��c�����>);��|��F�c��G�0͔z0�sl~=E��N�*���z��G��Mt��$$��eW��;ژ��t3�#XZU��xl�e?�gb��Ii78����i���}�O[�3Wz ˍ�PX�[��rʬ��DQ5&-�w�6��]�����T�ׂ������C�5�)I�k���s����A��Z��Y����g�q����B�}:���*�_i���S�k����s;A�Uf����o
�z�:�:WMV��Z2f4��F�/��!��
���P�}̩"���;QO�x�,:���}+���@�S�rD/y��L"��i�)@7
��(y @���0�@~2BT�!;eGgu��O?�sCȋ[A\��(?��t��3[�v@9����W�>JU��[��N�~K/�VGn���h$8�gh��>�_V�d��,�:=��2�����K��:�UjF�u�4��b�ڻ�J'4-=Fݾ�<aDY���w�h�1"�M��ӯ[���.Ѧ��D��cs�j#� �ė�F��ufS�*&V��AA���f��2�Km�f\k�a���ܞ2����|���!b�4�:;F�j�/X������a}��X�Ոk�},�)TP�\!��f_B֭�`?���6��S�3���0)�A�C����ƭ�ѽ{�7��=�M�J3f�Kh�sQ�\9��q>��qnL���Z�e��Z��vR�i[��	LFRjG�vK�kZt�<b���:�W���GU��J�ҫs����U��x��#�r��L�#±qx����案�����Hb�rk�#	q�zL.EQH���~h�=rs���k7�Z�P�c�8��0����D$�.<���
Da��n������,}���bR�~G!Æ'|Zb_��$�\F�6b����éT0P��WF�Q�on��5yT��[kx@S���8F�������.��ws:�F�X�)��!���b������ϖOB!�O��Z�t�����d�W�o�@5���Z�yt�J��Nju�Cq��V�*y���6���S+�q�Gy;�EI6�WY��]�H�[uNV�SH����G� kɾ�`c`��Z�K�7���_�~4����r�^b��}�����������:�/�x������Ei�=.v*5!.W?���8��*"�I�L=� ��R�$ P����Ta�%���TK|��$!S�;H��Ĭ��L'р?2�i�@� J�(�H�O���2B����:��ib�ɉ���Y�6� M�X��q��v���4���ú�;���m2�~�ӊ8բr��E�}� $��lTbW�w�5į�b?�t���د/ap8+u4�k9��K�7�\�EL�#�F*���FF��f��q0���:?*}��=��#��O��"B�(M��PvxX�R�[�0o�#X�s��J�v=���y�T�s���.%��v�np�o�!���Ó���
��M2��>�/�]�x���~�D����J_�]!فβR��D��\ؠϱ��Z�шx����(��Him	O	.Xz6�$������t0D4�1w�����SS�N�{Jh�KX����X v�ɱDO���w�"ׯ�f>?���-�*���I�Di��{�61]��I��֙i��������i�>VW�������E�/�A��U�K$,�ֶ��`��D=Ղ΂�ے��ە-<�X�������v,x�*2��P,ƹeA`�>�Gza�jJ��#��7֧�^��yg�\��:�Uy�ln43�h�@m����sd)p�l�%��t�>�L����h.�����fx-1&w�� @8l��?�qY��̽UE�4W�&��o�G�8	�i��N��U�!�)�"�y��(m9C�.%g���$G�Zi��Oƃ��Cj�#bٰO��l���k��;a3ő��͟7�BSn���;���(���d����Si��@����`��n"����rzjS�w�ش)�z?�z?�;��f��Rݢ��ͮ[�d���-�
1Qzo������tV�Nu!E�j-��K�֧�"���Z�b��y5'1���4�����c�ltVwp	*�ze|��O�T���!u;m��7a��l3�cU#P|i��V��H�y���7eA-�"�쌴��M���d+Ѯ� .s{�<�w3�"t���j(��x��*�ǩ?�1�;Tf���c�H��=�5fD�� k���o���˅��  `�]K��<��m>6������XcP�;�Nz#k,���Uj��c�-�L͖��Bb���+_��C�Jv����w(k�M��x���݆�l[է�6�� �������~+
��{q�ΒO8�l�G�P	��Y�� N�S�Q��kӮ�����	��iu���8��&�� 9�I��{(ZŚL��o����73��dySN��?�K��{�h=���M:�l:Tt�X�Ņ�f�<�#��UϛM]�
[a`������0�&��G��Y�ka^��m���K����",ЋG~��}����z�
��s��Q�����U`�*��}d����k�J>�m��N�!�taXz���TE,�W��峣��n�U+�F�Ƭ��s�Q�(�E����R?ź�����F�yc=�F�ē���o�����V�b��&,�y�%f/D���\����sfy�￩��f�ov��&M��e��&�fE�JN��1�������c��`%��.�{�R��A�u/a�$\��x]l�];6��1�kIAY�e�X���jG"���?d���V6hՙ���~�F�H*�t�����q����������c�B���[������,h5�z�&h�,�v� +Q�=ᇭ2��W�U/*��C���,��	�擊����߻��)��?�2���G'���v�0���yY��3J�`�3����w_D�S Ib;�_"?l<����P��o̰Mo%.A-��'F�GK���=D它���Dt���'���K�w8-�����M�I���NwC�����8+B��}�N�F�;:-�hj$:�n���q��id���8��+�EN���$����P�@��٠�9,�n(��T�eF�1a�,�[�sE��l��vb����	��Lc E��E���@e�-����3Ϋqg��u#�x��`�lr{��r.�LX}�)���I�?���ܳ���L�D`���lWp!W���)v�z��y���%4P3�l}%N��O���t�fwV&��U:��_�6W�%�K�v�qt����4���)a���~�gwM�r؁\qhXͽ�[�.P�/��05�:�6���r>�0T@P__J������J��w��X7� �������Ñ��LS�ɾ{ק(��|�ǌ�#{�ӷZ�����L/�EH��7���\R�o>��ɠ�$���d1�k8���C �)N�-�yE���gU�HR�,ZL��»�^�O{�;�NH�,���(;LT�s3�`�?)�����T��JB��{�%���š�~z�e��g��/7������d�t��4����R���fn��sxh$����!�
�9���?��ǿGփ�{�l�(ʼ^V,�3c8͌��$1��ܒ9,$րƶ����ȠK��9���=��,�:F�k8��¯[h�FAL�AmR�����X�e|��u?ej�����Ê�Zj���������ŏi�T�tZ�Eܯ'�ΐ2��X$�W�s���.���<X�ɂE���j'U��p�9�}�7�n2� �T�4��Y�� DVΝ�h�ȍ��c�=lj����g5>@�p|x�ҭ�gڛKvPK�V_�Y���U�Y���v�?�\���7򌴡c�
V���Y�?k^6��=k@�v"|�'���[X�f�Đ�FH�ih)�(;t����:;��!�VG}<�b8@0� ��	P��,� f�Fj�J���ڨO^T��P&��\�NG���r��_������_q�[�k���^IeVƩ�qJڇBqf�~�m�elB&��z�L�v���o�BV����Y�ܿD��w���.�x��f�F��؝ԏ���O��5[V�hR�p��w��M�,�".���4�?X�9o�ݬO��[i\f���ƑA�K��ܯY�<#V`��Dk�@@gJ.� ��Jk�������mн�)�tz5,Z\�`�ړG��VJCe��h}�T�����.NQ-���̶�������D���mP�#�>�4Ww�����<ژ�-8��p�Տ�#/����D�E���n}ǐ"��yw�^�rN�O�ckP�+/#:+!�v�K>���Ӓ�*T:�J��:sf�~0�Υ�.�\�(+��r���OK�:��q�8�g�$��̷(�>x�a̸�>�D(��
=}$�~_"s�짂�#��V����9[�аM휲5&�;����ȴ��4��oy&�Ƚ�C[���D�DĀy�i��tJ}}��������)�xr�M��~>;ޅ$�n���A8Q�D��4���<����Q�+��4An]�&�q#Y#�.X8�4�u��{�ZY2�[�y4�T��Ht��C����*8K��
n���7H�i p��cĊ~�ʋ0�&�L�� �Y�ymuQ�+�/�����|U=to��6��co�;U@���48�y!p��J�0��Kp����w�\Ca��?��`�+����գ������NS#l,����Ha��^�K��8C
؜�5�M��)���`g�Y��s������~4����&'�_���Y�q�6�e�Z�k!�xo*J.]ۿ�0��P�(G�
�\�Qi��)2P��˺-�Z�\�B���orQ.��������f�5����n���u�&5J���mWȿ����Ĺ�}Ν���	�-+v�\ў�ԗ��&~����I���y��/�Rrs�Ǐ�}d+�B�,�����$�	��=���k��ē�Ĵ\0-��B=��~��{n*szG!ꇡ���T�P���);`�r�������A3��oq4F#����� �m�;�A�7�)�~���FߺM_�k��+��}e��.ֵ��j���B�-��z�`6{}�`�M��pặ{��A�_[/�Y�����9=�?{	2S ���תs2Ѳ����F�BK�:��釜�?6��y��3"�V,h�ܫW���-{�`�(�ڗ#2.�Z\��v#I��]�9����G�Uw"���L_|�!1T�� �^����}����r�3���v�C�j煗9f �Cd�܉v� Tp���'�}���?!Z�RsZ�QF��zR��+Ps��s"+�:�鈻�A���Z/_��w���o-TF4]��2f�v�$���M5�ɮVY�|P6�$�I� �m$_]�u�&wz��&u+m9�p����O~p$&K���ſ��iS��*&�󁊑�O��)��s�'5��,�{��`,um����_�7;���1��A�fPٖ��������G#�5eK�Y��j��.J��k�'t�z5T�H:�Ǯ�R�p�_�"B~�;&��<a yR+V#m�p!�����B�r0����L���c�v��HE։iD9���'4R��<Ϲ!'��T��	D���M��`r{?��3X>_���3�i�}�g:����؟Z|�(���
��7ћoi1$�d$�Y��+���*���������6��m��_׸��s�7R�<�j-S��UI��z�����<����a��W@ˇ:#n:�.�]$�>K�G�d��K_�t����W�놊��O�Qb�q��]d���e��s����ЗJ��L�,���l��~ɸ�7���-]-љ�T�+�V��_ SR���4���{*��8^�Il�{���A�:HK]Nۃ.-�»�(fv�!�G�F�V�	D��t]D�Ŵ�t�ۺ���	����'A�Vd�29ӵhlq������&c
�\1�z����a 4a��a��]��V����\�V�p,���}�����A�_@U����:���*����G"J�OXW����xc�MKes�
�׫��n#� %O�d����7�n�~W�JB���`s�bj=�2߷|9��[�K����%N�V0�}�xb��쁐0��;:8N?˽���JS��OHdLٴԸ��E<���v���Ƙ��V�P�`�����"�7����<z��	^�}
I?�#. �>��w����Q�_M��
t�9���R��Ȱ��GS�<.W���g>�:����$�a��ɫ��6n0�.��	y��Y�`H�N��Ze��S�t,��'"�eM�@�����x�(=�@�'@�)�|x����&T|��g����tM��Xԣ�/
o�}����g�M :�]��K�Y��~�l���R��R�����sz>7�r�䄆�DPQ���D��lx�QT���>]�(�}��%]�t�t��	e�����;!��Ѷ�ԏ8�� ��W+S��hV��8X�`�Й���z 8#��	S������N����Y�!0>�#~s�>�hC�3KY�C+���n.�<��k.��;⒀(m�|]�T}�o��%��ɘ��4+��8������,�(7P$�>��Wd�y$�9��B�`	>Ԕ�rh��RҶU��R8�؜��~��mR�)��Pװ� �������z;O�[
uo�����4�	��V��[�{�QO��Ș�=L��pOKr�;7�D-�$�x&s�4�ć�./�)4�_M�=_�	R��A'��r�e�4JU'Ti�ؾ_=~����1Wq�w�3�������Q�4��ʉ#ߐ.��գ
�áY�p�S�8��JY6?}[��CG6�q�:K�p�5�-D�C�`��#y��oh!kD�q��أ(L����t��vK
�u֓���brcߊ)��-=srǀ���ղ�A��?�hr,��o\���2����.�|��Q I�	Q�6t��������#���� cbr�>� ���V���M&�,��$J�Ϯ��2���6���5�R��oC��2I1�D���iDfW��e�^Z�4/�&�:�:7?��=��9<Tf4��i!�u�у� �t�< 
-�>����CM�P����0{�����,�=�IIe�L1�@b��kJ�d``��w321��wL�]�(�p7�Yr��<
[F�D{1��[K7��7+l��.dk�����lU1��{�m����,MB���h����.����i��N���S0��U�D�Ez���崚�D����Er�qz��i/�HU;�_�U���y(kj��[��q�2QX��bM@1Z)f��g �
���YE�4c���Mx���D�xy��,��b¸��JaI�����}]q��Ր�{9E������k�g��oŧif��L�P/IN~vE��3r��k+�|ѿ��!��3ȑ,�Ϩ���p42�˒v}�Uw����+����s�a�dLwr�����r�4�e�qF���w�-������:mF��S߂�%���L(%��r�J|"cJ�_�R�����S�!$C�肼�d|���bD�~�Zj'8�����L8���쨐3�k��	R�i�H�K6�VD����<��a�g��,b��m�/1z]�l�r��-�x�����ħ�+����M�&���&��ΥQWd�����n4m�6�K��!Xk����H�j<X-}����S^����b�T��O�ؤ��x��x�EY�-��I�U�̻BXx��~�h��ҁ'���p��Q�߁7.�f,b����$m����������X�� :�&�o�ͶT�TZ�C�*�ypxl��OIcf�K=���	0�kB�Pr�#��Dt9�])J[w��Q��8�Ċ[�N,%��
@��A�5d��� �]��f5�����{^� �y�7u��m���k���K��s��_M[��G݂u��J�_����W<%�Ӆ3)�B��4��CC�QƋu�Q��/��#|��/�Idpwk檚�bz|�	%)�ClE<���CЏ]�L����M��Z��,��|�@����4�2Rۃ
�"�����$�RA�Kn@�����sT��|�(�q�����բ��w������K�ť�O{[����EW�Mr�2���uD�j��j�L]�Yh&�x���9r��B0wjsۅCҩ���a��3���'R�³΅��p�uy�E'ě�kX�������`�u�}���ie6c;(-�Ҧ/�6�"
[��h�)�\\]�?�ݒ�g�c���e��:&5��2����<(A��ߛ��k�+���@j�H�4B#���ځ3:bQ(�a�2�m�/�篟�ʸ���Wϗ=wR�v,���7f�����T�7,ڻ5r�'�<͠w�"(���,J���a����v���Q�K�Dw���U^I�ЃHü���'�����}���W�6X�x�)����.[+��	"w�=Ѝ\mx�0ʪ�!?�bf�����x�b}`���11k~�F3�hB9:��^���o��ɉ"�%.$M��K��\ًDsuh�n���ݵ��O��-�K�o�
7;-�����D��~�߆�ةEy���b%�7�2��{�������a���y�Dz�\�m�����gv��H��DXD�5�z�H��,H��&s��g^��j0m��ak�
X^��)|D'@3M����ۋw��~�v�v\�O~C������oJؘ�X}��W�PTyQ��?ї<�8=��}e]�^���q��9Q�$$щ����\H�W)b)�8�}!�����@}	��/,L�7T} W�Yզ����_�ST�ڑ�_�����D.�	�h(5�9�^4^�=����uX芋���|�O�@�df슍�^S7�WPB�@��cZZ�P�T9�<�����!�˄�փ��:�E,�z�!Q;�9X��.����=^R�;��*�ʜ1��7�m���.d�k�\���O���y$=n	\~���@�K=�!�
�u`��z�m�%ta��5�S����McW�I�=�b7DYW�G��ם �]`L��臇J� {H��&�V�,��Sd��c�[��B�`ؾ^g����$i�:�,F5�P&�}5<lܪ�!�����L
gD���"j4��Mp�k���=d-��>�$��3!n��Y=�*�9����Y�N����p�^��Ƌ	xH�
7�˺OuU��l"�	ێ_r��S�$X���Ƀ9�U8>�&S˰q���c\��6�F9���42v����O�����iޥ�.b"���lhe�O�F8�YR3#J�U[0����A�*hT>�^S��Eǥ[]-��r8����V���[&�G;��^��@�Q\�I�`�n�ʱ�+CD�{n4�2t�k����]qn��]�ffΌ���j	h4*nb��QV2��ۆ�����:�DX�V��f& ,�,���W/�t<^`��X��{0!������\k��0G}z՝����)�y���_J�xOq	�KW��So�<a�O�o�0\�}5���:.F���*{��[��9�!�s!(߂9/��[����E$�Ӣ'�GO�=�t����E�"���Ѱ�KO49 ���JB/`�Zbڗ��(���� <]C�ЩwOy)DnҾv�*p(D6BL�4(��ݼi:�m�q�:6�y��s����R�Ѥ]�d�r1�����M��m�v�ְ��}��(�R��l5t;���
�����pʵG���5g�OlՋ����46*��U#HP��m�o�r@���g��⯜DI4��=kp��s�I��a��z�7��ߥ��ї��w�@T��tx{؂����u��`S_\����٘��D��W�F`�nohz��{7�݆uی��+�,���Nb�j����N��χN��9\�mz6�֝~
�
?>��+�՗�K�8l	cym���o�#إ�EgQߍ��*h�I� �6��'�T6�}䳚������p4��<��"M��E��3��&��#�U�o��S�עvd���Ы�P#-C���?E/{�Lg�O)gGZ�jP
��g���}YY���|��%�)�u_��06��I��O3h*"��^���|��t=�{��a�nv�4�Vn�L��=�PY[ME���fng��mdgfu u�@�UFpZ'�@���Q:���k�}'��*�Q:k#�Ӻ't�7JXk��fcZr�-#�g��9ʗ�UbZ]T��φp�4�L"��w?��B���Db�2C����2��VA��;8Wc{{�v ���+]��9ϑ�*]� b�Wx��%��*}��#3�I�O���*��L���A��GWQ�t��]����9,z-lX�L�x����W�p]K�0%xB�G՛�-�1�I;Pe�~҉�I:��{tr��v�㿆�7��y̍Vl���"v>|�d9x�T���y�H
 ׎�q�� �`��`���*vD'��s�O�v_O!g%�*j)YFb��]���(���I�����ύ")ɯ���c\�Mz?(b��G�ܯGV`�N���2������P��䅠`�;���:�)�so���fy��@��IbNg±8�Kb�/�{��8���Zo(;�<��Ͷf\f��SV��Ӽ�1��t)[+	�4O���gE)�R�Vh]dk�B�}`����yɱ���c�V�����L��1�p�~��-���&fd=�G�`�s���W�h�M���* ~W���nnrY .d�P���獆&�]��)�nƫ9�#��gS�1��
�p���U������g&
������wTX~vBM�l�s��ӄ;b�a���Kx
���XQ?�=�R}�uಷ����Z����e{�|�;��y`�(��ŵL�*8&��}�<n~2�Dr���ڥ��l^������Hl�*����X�],�u=��F��%�ζ���t���*?��.Dk��s��N\����� 8!:��]��}�I��t�|��n��e�/"q��Y��4ɶ����^'���Y���?6�_C����hl�;��xS�@���>��u���`��l�������6�{���>7�v~k�`��4�9xN��}��{r�{!�${��@B�e���Q-�o���F:随�}���np
4�s�z���JtΦu�{F�&���kK��a���iu�����pC��Jқ���ȃ�Dd}��{����?΁���L���{7q�OKZ�ԗO�!l�9���˺���~�982�n�"�3'�`)l��ً#D�����v���_|��N���ԑ1��Ձ��ۃ>��F��9����-b]�g�D��[�I/)�-�&����=^+����^�X����4��C�|�B�d(��K^�j�%6�{�3-�-��`az������=�/�*���j[��Z��غ� )���giΌb��!AQ��qչ�����>6׭����8vY7qƌJ�����EbJ��7��Xt3�ޢ$��XOZὍӕ�i�� �����Bo���w�:AB��G�S3T����_�����Z�r?\�۬́;�ux�?��B���p,s䒞�i�
�ꮶt��B�����\���t���|QA��j��Ә(�Q�"�[�UT�}R��b	ݧ�����Ҁ������R�ʹ,�(������E���^`[y���OD��(����Ò��N�OC��ˬ�6�7�]S�A�3~�u^a�.؎���څ��8��/�����jA CD���߭h������89$�b(�����*)�����������f��j|�xE8�Z�q�b-]Q#gq�P����l=��F*]��g�(5hS�� ��������R��_`�c@�Di�U3�Hv�����xETd�S��hBզ��
5��l���| eCyE^b��"��܇��Kti��������Z�0�5�
D��Bvr��h�M�0��7�OcJ?��W��T��K��w��B�O�؄�'�7��_�o���s����Ţ�Q���*iw��v��ɳ�"'��=#^7!@��}���������j��R�!d3�n�A���s jGO���"0�+Me�wōF�`crn���;1��g���$�1W��zk�d !�B�u}�z�-r rR�Y�|���J$�"�8 �;�워$J7b�>(,�~G��o�uegh��I" ��RN�)��4+��4j�'�&o���:ٞm:�g�D���&�J"�Ć�����_�\\M`��!)�Ŭ,	���H��7�+����9~X5�-H�)�@34�ǵ�x��� �a���-��J�ud��2u"9����e�����vhjb�7J|��,"�	I|,.P>T��.���gl>!b�Ţ@��Η�A��HWy0�jru�l�X��D��\&鹺B�Z�uT�0g�A;�)�%w�o�2���D���c���k�����%s>f����-R�$�mZ�,��!*=e�����x*!�Q�7k#[��w������_�~��9e �AH�xpde�~��i���;�i������x?�=�Ҥ�
�sw��f�k�D���*�2��bH<�+�4��{���",B;%Ԧ�t���LTd�k�'DJ���jSffs�ߤ:�m��;Ǵ娰�zX��W�r�ǭN�?`�D01�-����IYօB@h�QCl�V�n���
��LTE>�u�T��x�֣�g<9S���\�-�E�H���ʙ*��!7�/jQ�"=�J�jܣ2|����vß��;��G0|�6Ip}��f�e ��6r��8�,R��랴�'��?]��������i�m}��bC2�[�Kާ��S�q������!���2�$������ͳI����G�G'?D�Z���/э���L^|�2�J��<⯅�n=Mp�g_<i�Q' 4w��9b��Q�0E����t%��ya)�8I��O�q��,o�J;aoN>8�y����C�6��I:@�ʴ=��������č���K� 2��v�_�rB�v���{F"h��*@��N��!ƮM���Y��Cؤ�������nc�]�War�>s���	�V�X%�&w�z,Ї@�-&�����g���)�BY���x
��b��כ�
����8lۼ�����>q"29��`�]ܸAz�|�%[į���YK9�o����v�e�"zNs��� :����	�8�4�'v���� ¿!�^�����e����I&�ӚX��u����h��Gmg� g̎o��yӭ��Z��xx��=e���HV}�s�$�i��p�������Ď�����B�#��e#R�EUަ@Zղ`�	��P4��Gy�� �JFU��L|��S�Gh�fo
�~y�GJn��_҈���03�t"�Hb*_,��Z�e]׊I�-�sӺ���5�u{x!u�	�"��r�P�Q���_��Q�#�Cْ��/��`�6�ޟ�~�����ԫ<NB�|���
QP��L��)lf���A�h�'"Ѭhw�.3U"9�:��=�?���k�k#��Y?��v���f<�raql�]�e�S��_Ϫ�	�:RS�E\Of�}�4�����Gݽ
l�	���ɀV�.P��ޜR�>d�_Z��A��+��l��o���@�_᷸��l�<�f"Cb�C��'��C����7�X�S���uK����m����e�Xk�=��s9�<��Es�/�$׀ �%�ML'���Sׯ<4䫑U�'v?�b�KWXC��x
�]pBXѹ�[a2%�O�7Z� �!�B:��tN���j�S����`�m�2e�jq��^mvt6�����J��##[V��F���	��.�K9ȭ��Q���#�XP`�3Aj��4�
��J��_~y�v<��������~./R/�O����?���sb�n3��7{������gT�X��o >����I���2���	U
��Ą�k�`�����WsH�����<�w� ʈ~v/v������k�b�5�t�`��њ��� �Jt �Y^�����QZ�(R�#*�ʢ'Ͼ�5^\'��1���'��WɎ�3��(d�yp�j��QKEc%��57�0�{��`E��l��i��`����%��o��Y$_� S�D�4*_��6��H��q���%�v�52�Lr�2�~���+Q1q������a7��瑜�EC�h����oV��΋ܼ�kp�`]?���";$r;��h�iZ0��9� ��5�"�G����i�c���#��-��O�G�3��e;���XO��͊����|��:��T��,o4�s'T�8�i�"�׍�_�(�������J�z 'ݍ�{�����=��%��&���C���EOK��i"4F�ݩz��ۍ䞝�<�GS�Y��N��e�<M32�C^��Bl986�D�St`s'i�����Z`ݎ��|�9�W���L�3"g�I��z�����n|���l�8��Y���I���Q2���`�Y��M��S"��OX-��.!��W�\F���SɧKlx���?���4t�Uu�����nd�V�>kA��`C�\�h��9���,Րt��^Ў�s�H%c�i|���5z��B�3lg��o��b�Dث-�|��Ju/{�k�c7�-'dv(��6���ԇ���~#V\H!�6��=�m"'�L-5��)���)y�V������������D��.㝸kTd�L|y�d��}���=����)����VH,ÏJ~���őt���@�}2n�)���E�1�wm)��L����%l�.��:���	G��D�N�	� ��]�_���%
��{�I ���Ij~̊��P���1 )FyTpЇ
f���ja�{�5x:n�)mL(�0����4�JՓe������Rq#������(��0�sr��i����	�k�~zq�qyI��_p9:uY���+��+F;>�;Э��t:�sa>𹻌�i���}G�4�طͭ3p12Wǀ��5n�E)G,r��s��ob����m��?r0g;��JsO�k=4���-��;�{m�t�������3�^��K܀~U��Q���Yex؊yh6tu�z��T�W�h��=��\����UK�V�Dtr�h����)sK�*�I=L��`���ck�_���z� fVyn����OQ���g��5�y�:��j`�a8�ݚy��TW����7�P:y�a̽{'i���L����^���?��W<N�?5B]���0�ͯ`�������f9��^��h�po�"�&dS�@u�D(��\�+��|_%y�?'y�f�3��>աn=���I�O�.3�	Q�&-z(h<0Mm4"_̾*��8���!��!�Z}�����R �؂�X�(���F&�����c�3V ҈��������Rںk:&�d{ng2��X��pZx Կ7���4�=�:>����=�z�h���aBȉs�"�)<q��%���\I`������3D�����]c�Z0F����f��\n�nqΚ��Z4���r�luD��@%j�����_5	5���%�Y2/5��i�H9���M�d���2_Z�,�����~戆�����Z�J��V�j܋����e��h�D=���ctg�@�h�e(dY6����v�z��ċ�"����=�tp?�-/qDV�RhC��=�G��D�cᛇB���9nd?���L+zB�ݚ���'���|���Z@�En|��~�=GSa�"WYO����H̢��r�8r�����tVu��C�9G�F��ۖ��jD��e����o�[��v�t(�ݝ����̅�F�#��Y
|YBsn��@+O��$�5��I��r�0����uH��>)�[�͸�'��u���@%:o����gY@-�)�j�����؎W5�
��J��}q`�h�9As�2�S<���A�FB�_�a<�
�I�����<���Y�ُ�&�I��n~*�2��+�,�3��(K�D�~"���l��Y���J�j"�����U���q��V�䨿��B��;|�Ǣ�����I-�zⰢ�!t��&��P ��a�qB!	�7��k@�G�J:����qf�����IV	����\�O�T��/��-nn1���L)uU����23��`��Е8X�Uն�@��G_S��l���N��_�Ê�Щp����h- O����g��&yLz;��(�b%����.XqJ� �y��6'
��"��9	�⚉"C4��-k��7�-���(�[���KW#�����lc��lK7&W�?X%�9�@���6U	��x&�Y�D|X����}�ͦ:�0T��b�p}��z/��t��`O6Ye��~QBC�nk���<�jg����f��I4s�֋{��Ҹ䢿f�;\��_�u���JA��x�����C�y� G��L�&������0���*3�N�/([�����Jg!w�)+2�K��d
t{��G�3h��t��=4n/wJ��iW�B���6S�'�Tp��`y�G/qDI����1~U�w�1ܼ�4�������y��1vy��㓷~�� �U �䄌+9��.	����9���@�C�FR���<���C�[�p�|e��O(�0��(�^�3�1<>ze���b�a��@~��O�������_��܋�Z�?��$x��5�I@����A���4�<��o��oN�GWjfNc�U��瓼]��1��,
���O����zπ�}�31�C��'fc�.��1՝[V= �?�j��<yi�A^���@�3>Y��a����(�e4,*����x�=����*'�v�?��J!$��� ��}��������{��pk�	�u)콈K6�S ���&�_���������J8M���}�;_:�}N����[��vו�Š�n���#;��.�d#['�Ԇj3�~��*���e�����$J�,K�[��Y�eV棺M ,	V�4��T$YA�7ᙞ5�E ���6��3D����&:ՙҏ���J��^HqB�8:")��t�d�$-"(��g��O[���V��n�̬��- ke"�AW�*�DԲ{9��IZ��q�}2�ew�Qؕ��#�*��$�8��{;;��nY���__ˈ��a�
�&�����������Y������<  )���]�U���8��CB�?nO��.���}I��Q��5e�W��f@v{D�z~65�������XΙ=ӏ��Ղ���6՚罄6Y����jT�eǔ}�_��� �Cۅ mj$`ή�����D�l�Y"k�O��ܼ��=�B�W)���I�Q��J�0���@:�C��i%�ģ��bo(\*�Ty�=bJ�#i�����+��`��b����9��s�@�)���K����H�t��j�8y{Y��(��|�aog��!�t�p�L�a�HvE���>kl�K�S�c�OX,b,@����<����)vڒ�ӣb֔/�����q�Ʀ�:#�49���%��77x;_�b�+@]S�L1���`��#���X�-�>��Փ{��r[]y#ҹ=I����&*K6%��r�|�HO�c��kx07���Q��#���h���MBlxX̤�X����Aeޙ���).�HU�8hCd���۝V=��������U����X�+�-��Z9
Q��F��T'�;H�A�W���8��[
`��V����𿰿��,!�&����Y�ٕ��e�">��Y�~)���.5�˔J�<.,�W�VG�ה*��	1�Q"���.KeL�U�w@dZ'�>ꅙJT�x�TE�L���̹��mpTg��@�:��=�b*8��l��~p����i0�]��u��J�v���&#������w:��o`������T������ʤ�7_���n�Ƃ{�{u�C�V��c���F(2�:@N�Y��:�Y)�"Y$E�_g_%�#�%��[҃�{�[_y�'�u�	)%�1(2�1��k[���8���R:>{���GfK��C:�>/�	W����"==��TE�)�� 1FONJ��lz_[c���6��D5��p���Ȩ�M%�^ΥhV	��Ӥk&산0ա��x�ar��h���I�J+�U l7�Ɏ���2��^Liu7��R-l��U+�eQ�,7댾�¨� �cy�t �ʫ�wp��*&�⟤�(�oa�|]�'�M����a��Xa��A�~霿ڰ����a�
we;�gs9��L�8�Mw��p�II6�G��G<$�HSWƵ�|����h6<vJ�N���Kxw毐������7���.T�Ԫ�����n��^R+��uf�uC�d*�Oޒ�s�}C���6u]�V�^���V����'F-����v������D܋;��۴�o�Lݶo>�_@6zL�mWC�=��]�L�����ǂⷔ����&�o���K�we��<n������wϰ���q���]X�ߘ��Ey�;ރB�^��F����x�q�A������-܄�A%ܭ�w�����.���ܵ��ct��������L� +���L�4Yn{��\qI�ö�I˿ �)IO����]xre����
HV��.e���7d!���&!m��D/�����Ӵ���yP����	R��:�-4�e��H&wl�L�h�t�	3Oi=7�xE�i�T5���'=WT\Q�n�^��z㥆�!�v3�$�\�hU�I�iM�'7!�����f�\�cۅt���OO���B�b����.R�9O�A괦����\MN��6���0�҇M���zj8�I�Y�1޳7���IWm�(j�f��
@h:��OiKQ5�#A�8�DhP�RN������elہ�N�z�p�����:b�h=(4�9KDem�V$c�`�z����K..�$�&NR�+�3�D��M����A��^�"�:.<���k�	.%�}�Ș%urn��g�:"'D"/g���;e���C�N�$��D�1�~>P<��H�:�tcѳ�#�.^��n��Dv��j��V���'�\v~�����v�D���8u��l���Sd�B$�Sڦ�SQ�ñ}��sY�KL-��8��V�A������غ�%������E�������݉A�
����<�8�th�Y�^]<����������pu�0{��oPr��JLD�S~�緫.O��o�(�i*�t4��ǜn{U�B�T�t� e���D;H����q�R4)��6
=�k];�1��ǈ�| �usP��5�	j�D$6�G�_�}��Qf=bz�/k�	�.�� ĉ����;��G
�A3G!@�ϥ�D�bi��ܿw�V�1�R�4��=wb9c�eԊ��K��{��yVJ�,�aς<$n��E�"��}�L0�����<�ދ3�,Pe.QuAw����`X��Ռ�FԪ>7
�ڎ1�0e-*�BZ

�/yż������ӗ�n�k�����{tE'����0&�߁`VL��x3���# c<���e�MI����w�A2d2�J��y��P��.�[��wY�9UH��'�U3�ٛ@�-i�	[k�I5f�[�$sz$`�24L��ﳒ[o��m�A��/��`��\��t~�q��f�T���(�б%�F\��r�A��1��a�`���-A�]3<���}G���o�2����5��Tv2C�豑��.��< e��<n����	���1�&�aPG�H��"��T���g��ш�=\���
��렗!|�-��������Og�䗦,"��z0�����Y�d&�/1T��)��-��	���V�u���*�^�j
	GhV�<�PǊ������K��F~�w�5��I�K,���� �G� �p�.[{�=M����dK@p��,�� !p���r}�#��ϬR)�hs � ^�U�N {���Gh�LAE%�Qև��;V0��t�5:)H;>�����'�_����;��c�]�}�z��ŊL��p�''?�nq��f)���!��jM�}B�n��l@�<x�Pӷ��w�Dp�eUh����
�>c9
��A�J������.��u�2e�cEO�r��Aue��H�,2}�����!|�,�7Ѿ\��2��/�1*��c�?>=|�u7�6Y:QٴQ�>�5E��>�T_�/�N�)YHt�u�����<��N]�/n����.\�$�
�v�ۤ8M�.����̓fs�$mg7hU���#v�'5�P����1i��G�%O8��6��i�q��"��B�p�2Ua�Q�c���p����`A������R?�85���V������@�.�)#6Q\&Dv�0^5�¯&�j硪Pս$t�3B:}-�=��u��`��L�N���B"sQx�&�SI�H�h���U޶��z��A�21$�mfx�t@0�O<^�	.�
b����uyl����5F#�F]�����A����uo��&n��R|j��q�k{}ˉA/c��z���<�iʶ��A�AӨந�~���
	�� ���yih�5��w���gΨ��dv0�z��Ї�8���;�C&ߝ@Y�����`��jN2�o\;�B���o��0/?�������UM�Mk�+8��o7�其,���a��m]�e���G��خ��V��j;���R�aF����~� )�8�������{��և��j'�N���ٲ�;��H����8ٴ���w9�_J�P�Y�.h,�ңN�_3衅p�E���)4�IDǩH��Yfd���)XR�(�|�1�_�VS6q8�E�"�7���G4�xAb|�EOa6�'��RoB�IT��cm2|���7Jf�j�3��߀���:��A�����)�I�ҹ��`�nL9.�"�-4i��R������q��X�a����l3��B�Z��}Ӣ�h]��/�v���}̙-���**n���Sq�-ѩ��_�����׺v����m7{.���\0�zX�e׸�ﯢ�`��"�rJq_�� ^#m��	r�>���IZ%���Ej][dj��j�X�{2.�S�V�V?�t3��	к����:��!�"� Y;��4�F�Q�T�@�8,
��'EK��+�%(��'	���\Vf!��|Φ�l5e�;4q��{΅���Ӭ��.�;a�����ud1�&f:bd [��-y����BT^$�<����:J��ߢ}[9+=����#��j�U��gst��2�RQQ��s�XY����*�>s5���ޫ	�(�����kC�@g�ϔ���8ŵS{Y��d�?(�mf���Ă� �^�OD�ޫ��z�5Y�����,�9IW�x�0t�{�7�f (�E�:����i<m�LX�྽�Z����D��k�\�#�%O���������=W|2�>��?��8�0m<��	\�;�}/�7���a��.��M"�,������l�yMT(�	��[�ۂ'�M��S�=�f����W,�j��aaM�/��O�QQ̷(��ȥ3��)è�[F��[�Q$��qT�����R%g������]���bރ�����v�+��	 Y��ٚ��2_�
:����y��Ǳ��
�f����cElZIi>G�=�i�������e�yΐ�g�Q}t:�r~��3�����i�7]��*�8bV�
�*;�o	��Z6�c�)J+^�8���A��RU��y�I��Q�"ƕ��rH���$c�c�=Wp���]�M��,,�� �-B��Q����H0�Ƈ�|�/4A�=�?�|��әtPB�NQ�䙲��\�|�J����Ezμd_a�j���7��ek���~_+���=�L���~��g.	��&�4�q:��w�6���R������=���f:�v����L��@w��pGY��5����OG�6�FޫƼ���M�=��3޽$Q4��X1>���{ �i[(H
Ap�s !�nG�9X���k�mvA����ƾWg���gX~��'!3"���c��(ϳ�^t���5\��|m�X����� D%�'ﭖ=�u�� �l����#R� �x�ӿ- /��x���9�%_.��wI����o]b�5��գ��^T���0=�'���d1 �4����
�|.���6����rmx��Y��LT���N� �O�ߟ����U��8ꗛ���9/q�K�����f��\}�=�4�1��e���A��ޜW�'��	2��k�e|��)�I����ڠc��V��v�	��|�b�J�����HG&&��m.��Lj3�X8Y�e8)���}6�4���HW� `Z���B�����V�J�w쵮ɪ�A3�汔��+e�Yh��+?c��
=!��UJ|�y�=W�辭m� �Y1k�
��,�kr���!��:�l�E���ޭ6j}���9��k�3I[&�)ʊ.�˞즈Sy�������j�k��X�h^��;72"`mU�?p��q�OcG'��$��h,����o�?���{�O�I�3-Ӕ%��ǥ��#%Lb�=^E�`[�xt`��Y�x^�����(��_s� �Q9���N�S��)�|�i���e�&Ҝ��	�C�������H�jg[4��f?�-sIo
�xB�Vu�s�|(z�LS�յ+mp�_sZ�aǽa�^7Thg3��Y�.쇭����ـ�=�/���+|���L-��GP�0.���',q��Nb���H�G�~�p=F��3�m$v
E�����)m��薺e~����9�0������}3�CC��Ѧ@�Et#~��i�;� 㺥dŕL�[��O���#�����.(�C `�����֮�M�N�D�娃���#����f�{��x��CH��y	zv-� �L�I SSE�pR�$�̗렟5�r�ެڏ�
t	.��R�����ጣ9����'J$iR�u�ς�oS���N/yS2AI��1\$n�3��~h�9+�G[��������Y:��l��A8*�X� ��z'�.?���8�Q7�v��B��S� �e��4�՚K��jB*�]��?�In�͋�ؗ!D�{蔉���IH�P���2sݧg�(e�[���_���t����"N��J��(���Ū������m~��N���ہ|7��/�Ư�r�B�">�0!H;�_�c��(��6� ]�$iz�b]d�;�{^*eE���,*��#*Σ?+d���&�l�ʹ�w޹c�ƅ�<��M�ƇǉPR1�Kw(��T����~���7�J��y�\�&�Y�c��g΍FK�Ǡw�?��E�ť��g�#9�_��ѢM�	�2�f}�����E��h�je�w���ꧮOň��l�T�p�o�2	����*��7yޅ?q67�"���=gxڈ7�Q=�U�E,���頙��X�����(�$�1��_k 	�U��=!���Wƍm�r�,�`�p�?f{}Z��� ��^c���O�ˎ����$H�����R��=W/nu#V�?Q�i�O��$�`j��QC�y1LĲ�ʏ�:���%��2��� r����6)6�-)ު����!5���[�W��=��1>��*8�� Uj:��L⥚7xN��\��zQ���b�e��˓k��U���.$�}s8��(�Y\�I��c/`� �ښ(#r�gg�3uML��t�3��2az���%5�gR��qoe�
qǶ�~����@���	����;�}���@�X8�Q�@ּ�ql{��n� e#|��U  *��ΎK�J��RYă�� zzs�25{���'�m�����7Fĳz��H4R���'�(d
k]���J����Mh�,��xKQ(�q8X���Cl2�.6�Q�5��a�����z�ǒ�R-Œ��P555��/Ͱ[ʢĭ��/�pl,��,b��A��Zo��2xi�0ЀM�M�-���f(/�:
�)`b�p��<����/�f��39i�?��u|�+ڐ�)�᝶�2T-vDK��֯�����Nq!^�e_ _�ܛmƋbDb���
�6���aN�s���ii��}���������Q6g6F	�uu$�Q!ta��ڃ�<�����Y��|tb#�]��.��qn�w�np����sOA�mnݿ���h�K�	��`A.^D�Q~�L���Y�zI�(���+OP��ut~�.m��Ų���u��T	e����s��z�?�~h9;A�1�y+Ƒ�育���"���*��w�1	�����ք�k��^����
��J�1
>�	�P�?l:Nhh4U�P�q*Ⰹ�;X4.�����4&�D��Kp�Ys�2�3;��!:	͋��������^�R���,�q�����w�|x{�h�=A��I̐C��뽐Q8�t�]u��+��p����y�ѝV��˃���F��EXc�>�����^��:��ȶ%J@��S-�{P {7�D1��]YMuo��Ɠ����¼�E��)n<Z}_�!:���U;�w��j��S�Bl�t g>�u9B������{Ih�Y�d[�xFz��Ke;��lQٻ���.?�ڗ��4o���9���CD� ��7ŰDX��3*�� �h�4��c�ND��	��m���i�����ߣiUѩ0f}P��J~��Ũ��}�Mmn̠���Էũ��_���(�X�\���c_�T��f	 ��k��О�~��>�3$Z��U z��W]��@w���U9�����w=��%Fpo�ٸ26��l#��(_T��UT�&/�5�H݅IeJ��ZNe���9�Q�C��E);<�<,��c���� �עE\Id�?�!�֡�!A�������?1%�hL�Ԏ1SX��fS��w*�l�)�"�/O!�$��?ył+��ħ+В��(��_��7r��h�q��g���A1�V���ؼ-�$���~���jn���Y���I�^�(Hy�`թ���q.m��Q3����^�������4��2�Ol�Χɳ���7�8{%����Ks�Ĥ�T+����ڇ��3��y��~��5w����!��Z2�,D�O���NY�5��_v�ߞ�I�k>��2A���t$ !+�FcBC-n��y'�h�I��g��wM�������0?~�x�����8��]�	o�e�h|��V�|�IZY���ﮞ���c$z�����s/�U�ry�E�3��)7N�_����;����K��׳ۦ� ���Q\��[�a��6�BP׵�x�3li*ߤ��ࡾ1�J_,]w	���婟��IN��ߔ3!���}R��S}Z��B�$���<~�$h���M�o���9�Q�T�i�j�χ-�<N�%�P�s�X�qY
)6KkO�`I���UoG���[��ކx�MKI�	~;lE9t'd�����d޹�S�z����p�<�`��{2�'p>����=r)�V>9�~��39��4���� M�R�������*���^+o���o)���p���ҹ��	��<9YKU��Q�Dc��9F޼�nt&��f�TD�ٱ�W�LnW���yu%Kh��Ė��|�o	�/p�:�1U	���^�����L���&��k^���ή�yRwm��tl���k]������`�a�,/��H�[�DQ������l.��Z����W+w���M	;?E,e����'��ϵp�z�+eM�]B�*S��d�찰@��]lc����I�j���2���Ⱦ��	�+M��J�`q�������6e\����M'�W��Z}�K��K��c$N��^H�M�Y�t~�b�&���3Y��?�����2��t��k�<C�r�������"�cO��Ή�yE�Pu�j�n�G�7�|.w��� ��J9���������^@���p�ύ�<��r�g����>��(l�6����L*5I�2|P��7{��g����(��\
ҷ作����XE|���Jv�����_E��HEѫ�rξ����R�mbB�䲷�9�ݚ �5�x%-��}��[��Xa]��`!Л���̈́ޚ��nZ���'��9�GU�83~�'�th"�05�.	~Z��L��̈ك��v��ɋ_
_�g�(g��߰s�l�6�p��_Sv�H���MsWJ^�[/�/��� E�dLp��?*����$U��^Ԑ]�j�\}ET�C���&v��%�(7Y�Ө7*@��죸c=�dO-����f����J�/t�4�#�0{a��I�5Pcn��$5O�T�:�4�ErJ�|��t�|�j_�\��?f��-��pV��7��s��e�{_�q�A���r�Z&$�V����f|'QP��,+JH5%�LB�
�?5�UI�Y l��[�nV��܎�r��Vp��9���ݲ�Qw�S
�=ʸ���S�i�1Py��գe�a����k�PM�˖H��7,'#�A���+j��\c2�����EES�?����\�3[c�0�):i�q>�\���N�]�bSa�{��`�!m{K��Sb|-����j�@NÈ,�o�M�&�gB�e�|����C�$Z��QF&�����*��U<�k�X�t�J.����S�X<�Y��pfd� �YT�����y�Ϲ,�	db�W@� �؝T�Y�Pn� ��I��_���X_�h����8�������I�I��ƴ��&�+b�J��|�Qh�n�Q�Ӆ�k'����M��X��OV��bP�z��=ȰpI�-��X�'k~&�Є�UښJ
q��l�2�&a��E(�q9w˒tJ?���	���Xvr_�1�%�=+�����UMB�����O+ڬY��o������~�9����s����$=�@�0�Z��%�i&˃6��^�8��7� ��a�P/Oh����7&�-��);���~&�?� ��EV�̰Qم��t,�����ਮ�r�N]�kV��Y\�� ���s�D݄�����u`A�]f������� ��p"0;��c���h�|����6��C��pC�׿��Jξ�Xt-�M%��ƍ�r��\xRztI��@�	1��/@�t��$��k�����Oe���6���
h�<�!EeP����8�]v�1��`wĎ���U8c�>�
���|V�'�|�vy#}��b���|�r�PkƂɎ��p�@���JG���ڲ'��Kh@:�p�3���c�|�X�2Ci0k#
�~o��SѺ����N������^���uzLv�M_���G��mF+��qHa��V����n�73�:   �.�(��T�Z=��G�����p˃���kTe[uLpB�)�|�H��~���~X}������^�h��
�������ēQ��]���L6xJ��[̚�9Z*�� �|����w��っ�@?Rj����g�`���,�
재���K�}��qHi�\�������#����,9�6�PR�����Ѧ_�L��~��i��T�,@	*� V��(�Dfy�LEl[E�F�.��_����4�]�c��[cmqB�L������;��Db
����@	�mYv`��
>�K�=���V@1��ie���XV�fng�Uב������H@{e��p��������fyh�$�\����_,>c�� lҴ�=c�ϸw/�(���ب�Ru?T�e��d�qd�	Iz|X�:���k�.:K��� p�zR�O�u^��W���m���߉����?��Kd/r��܀�����|W�a/�M��:[#ȅe`&�@X��{�Ô�/}}�%	��˔�]v�5��
UVm��/0�r6dzj�?�]Xw����,B�$���6uK9��3!Ɨ��eI���3;�ڼa�<����)ۧ�7᪢į�ū�'C/�pi�H��{#h�>�H�dk
[43c<�z@��x��b�#�B�g����W'�>�Pw�W0 /��Z ni��>&�w�����w��n$w��eMPƴJ��Sb�k�حZ�r�>2�6F�L�@Sm��;�?.`�V�P��F+�YG�_Y��\,��GZ�����xp�"�U�Ŕ����j���P��귺T%Ƈ�K�|�t���	QZ�!6G���!�pq�K!;�yZ�oy�J�1��v"�[5F��\�i�b`��:��a��[GD0�:���[��q�Ry��[`��X��+��wx�����8���Y� Ү�r^�M�ѣe+�N@�p�����Vx $*���CQ<�D�s*� �ď���R�e��/�q�[��mX.���}3L�6�1:�G��[A�2N�ؓ#�ȋ$�5��E�Z	U<��gC�Ҿr��=�$��/K�� ��b����{��x�Baz^��
���ZM�_�m|�������/{���ЫM���*��4�Ez8~��˔gQ��;>�TIh�W�M�1h�ڨ-�m�10��5(��m���T8�e�CA��m�����g�r���s�Tk�&`��$s�łߝ ���%g�$��DYb,����lU��Y,�v��=�a̹�o0� �����A��a1��ҋSޗ;���F	*c�&�����T��`�%H�C8�K�޾5�˲0�J�C�K4vy������E�,{o��
�T�����Y�_Am�,2t�����hn��/!J�x�։�8�B11�,!_3{��ps+R��,O��U2&�y�cq����YCb�O؝�!���;E�A�!0�6+�ro+�А���ګΊ������q9~�Nq�c�a�6�k���Ϥ�=��9wXKl��ځ9ה{c2A���7��=PH����)O����Ps��b��di2&q4�:{U&��l��"�V�`�$ڠD�R��R��$��c��
�E�Q�TC�q`C��u=-�k�į���mڐ�e�t&X�3Eq��%���Fd��e���W���"+��щ.���V#��8P�b��J�g��`(�څ�����߇��Z8� ��(�}v�T��;/=�W'G�T d�<p��t\gG�:�2�D}��$�߽F΋ɜ����)m�[֙������ݺK���y��o���#�zIJ �ҹ�hVّ��"b:|Za(��UE�,�q��5T��3iw�@��	�P�4�I7�C�\��R>����tO �ͬ��|La�1��Ss'� �:dH�H��qD�PC��ժI�z�x����K���>��3�>�%\�C��y���fJ���+���5(]N����e���B�T'p�,�C�n0]ӄ�3�S"�fh	�	54�2���9Xz�l�̚��D��x�tܖ�q}�-�N�l�FL�d"1µ�'��2�ϣ����-�����,2������/���ۘ�J[��hpȉ}ɖP�ǐ\m����w�9 	��"��w���O4���
�z��L�rW}���f��H�b���%c_���^�7^�ka����W&�X�������@R���)=P={�=X�<��o�A�e�+5��s�{4,��Hˋq��fQ�H�`lZ&�+Ђ�wWk�Nj;
@Gn�
IK�� �rQ��简:"��K)lɆ����hfK���$I�9V7o�p�2#B�>�q`f��@\���L����'`���
��B���pW��N��U|�o��ߢd�`�RnE4Ӂ�����ߩ�pJ��<��x9>}�b޹H%Xp�9�ځ���v���v��T���@�i}�m�;D^	�M�Z�`)���P�9[���o��#�/ԩ.G��wZ���9��x(�qS/�4�W�'#c?��E��/��'%��P��R#6��!ѧn3�#���g�υ�r.;f#�`�����_�p�J�H9����jmܼ��I�/�������ĉ�W���`�ⷹ����y���	kW�:���'��W�)+��
�u�%"��*���
ԃ[�n�E��$�ߚG��UzYn��ŏ!��?gd�w�pa��U{��W���J��:�Jv����w�:��~����ar�;�8��B����uјb�N"D�}�o�J�gէ昆g�P��k��q{:�E���+w7�)`�b' ^�].q�U�2��P|���� ��~�,�����!����u��4�q�~ɍH�%
�#q�Ŏ���&�
=�+��We�@��?@V�!�H�y�|���S:��'��U�T��<�<L>�Ru�x��6GZ/U�.�T&.cY�Hڅ�
�,!X������Ti3rq�����G?)�:I�wE(E��P��r��a�oO�!&O(*�k��,8��!��!H��� 1Nx	j�\��h�b��C`͛."���g��_�Ƿۋ,�|�J|��˺[���tg�U���i�1n���	4�8�'�ϛ#��?��Mn ��̭�s��v�<x���C�'�T ��y��^���MW���ޢ�d�? �kr$Sb��̖S�`_����E,���V:a�KY���U�|X!hwp��2��/�D~kԘE����u��d��U�ZUN!ҕ�{��?�??�����xt�6lKt����9��b�m�#������yJ	���ՆrH��1��[�.T��q�Yt]	�O`i��:�΃'^sZ���5��xCuB�){�ȻO~�<�Q��ʜ�.ܑ�3A	�����f��E��e'�]�-<���Y"�9s� ��u��Κ��0~YYV�]��yA��a&-^�w/C��S�h�7�ٮ��f�b EYM�Kn��Y� �i��+�Un](�c��n���ꛈT�CIK���x�a�"�(�B2\.jQ|� #ru]�B.ಏm�����4�䎙���H��u�����'X?��E�$Ԁc49��:�MU�`�� 1�2}v�^�7�Ćh�{q ܸ����| �*J5��g�9 6�� ����ۖ����f�
'A�nT���H�sv}/�g�����e�j��bt��|[�$��l��e�3oYT��بr�94x3Tlw��z3��^�	��&D,�
!�� �,�3�2W�"�෽W}gB2reK5�헥&�R.�hh���>rD����V�J��CnVg4�`�L}uY�2 1yFO�/h��I��P>��}Hmq���3����Dn���ґ�+n0�\���E�q$�R|ᚓ�H����������!rW��/$a��Vp�����}ɽץϛ���ft�����pY۲7ƁS�޴�0;�D�5��d�&t`RaJ-���fՙ[VQS�F����9������M�f��=��u�B�K��gw�k:�BJ����ɠ��=�<xaA��{� F���R��ɘ���	8�'J�U�ۦ����r8F��=r���pV�Q�tk6�����ԅ�E{j����ӏ���XB�%- VB&1�*�s�X֝��ȣQ�G2z�ε�/��Y� e�	�L\��6��z�3-�u&�M��	�0����dz�hߩÕ	U��~4�\{/S�g��b�ew��~��ѯ3� �qc�j��r:3�:;�!��Vɮ[�d��$�~���Ŧ+�=<��������d�����Z�]���v��U���Ur��M��ǒL�<�["�^~c�맚�S�ӷu���>�l�9�R���rJ��v�1�z_[��ɔnﰧ���߲���@c3(⒆��0��D������.&�_2�4@�\zRX����6�+2R����vOlO儷*�M
�៽�� bY���i��l�����t���3��IV	腿J�mp�Gܴa�M��ȥ?�=���\�j��M���ݽ٫�!ʧ3�j~����%�S+�#�,��ǧ��4��ݸԞw"���
�Q��;8��lV��n��P�c��t	��iy�!�,�4�
�Aؔ�"-��be���3�b^'G���S$��U>1�����t
�=��A��pQGx����Yo��h�r�Hen�L3r��gD,��[S��G7m�.	��+ɕO;J������O�/|�!p�:v�}B����B$��S1��"���{�x���m����c��2�j�\�7��i�:/�i��2�W��P=�`M�	��w���3�`����7+|]C��I"5Nɿl>-v�p����KuK �U�<>Ob����ǣ6l ����9��Z��&&bn'"��� �K�J'y"��1�����8L�6���S jl(�+�*�x�6�t� w���	A+C$8�~��h)}�4���N��v$���xN�
�/���֪�=���ǲ�ې�� $�5�p�M�c/�d���v�*�?���y`��� T7-�_�tq8V���1>�x�+~�e
�q�:�g1c�J6R�����Т�ߑ�G����]�tnlׂ�����o�YI�2�C]��DA��tb�i��͎=��ZD4�1��rP����s���z~�c���V�Y��rR�X�!����^�=@�ՙ�f�ȗ��θ:C�Ņ�s�+65����2h�̋��f�σ��n&h�������!Aų���1��ôPȊ��:����j��kN$��T�&��4?�S 9�I�V�UYs�hD��*!����ބ����)<�j�dI�������:�P��V9�������I{G��s8⨐!J�g/6��/� 㶨��B\� �n��!���F�t�_�T�D5�!*�1D���e��b����C�
V�M7B��t�����#N�C���l[~�����Lxvl�_��a�z�'��X�-�H��,0��a�������,�Y܄��<�HX��.#_iI���� 	�� ��B �f̰e�����-f*A^��||�X$3q�SQ�����
�L�S*m�<�@oi�,U�Ց�_9�d~u�?xh��j�m7"����Ob:i�n�����A�ښ�=������%��ZS5�Lw��n��X0�/EqdqU�C��v!O�Ļߨ;�L@l�z�{x_N�ñ3%�[�O�|��M�K?j�(��m�0�;���MW0̡��/��Kv$Q��t����U5R���;y@#��0(���-�K�}�S)=��������))F(���9����Q	���f�;���\��u+p;*5���,9Ċxe����+_<�;IP��m�7Kb���v��A?A9x�t9iM.�� t��5jZڄ
��ݐ�yXu�@�}uo�F6/�z���RM��Nu�5�2j�����&KQ���-ر�Ѯ��4�2 �؈K�9��[�~�~"ҩ'���@�-�7C���!kE7��l���-lD9�̝�9���}�k�^Tx�C(N�қ��񖭤$/���3
�aWa���M� #d-~�d��fٯt�"����=B1�W��g�8��_qO�9�a�WVȰc�ˍ��aq����7��=�JCW�����D�f�"�gG,?ݧ�׫��tI��0�K1�X>������2'�*�$�K��������콯LD��ʍ�Ԑ��p��x�qP����*��� �1E*HHv=p�7��S�s8�9�xT�А�J�� 0�G��A�<�F>��i"Cܻ+��Pjf_��dԔe�s��h�`/E���J[v# g�)�[)5�Z�h{yd�B����ᜳ��l*�-��йQHT�`��cjo���D�~�k���������e+����'��X^1��GK,#���[�.�?��Q;�⑜��^�p074���>�=�~�i��$�LH�5�R^j���RQSRt����x�eL��]�����2T�������܆ՃM�I`w�CS8�h&�;���!�m�Pz	P�TZ���Dl�Z�o�$����T�c[�����_>E�~�?.j�p��?)�M�wU��P <��.-2��w�$7��P�).oSt�Fp
g��F��>#?�n��;_��`�o�)JZz��w�;�į�S���������%��2l�F��s��Y����;*�g$�7���0gsO�����3l�z��{a,��;ڊP|��iGj�%C(��c:�ώ�E�W�)h���W���KJP�W�Բ�$�y�N߯O(���,�W_�)Ity	�gmI�x��F�8���d�k/�q����=��,R��bo�T����d]���'��|�"diC�Y�"�� @@{�Ԝ��
��18rǼ��}0�	�~�V��wKt@wb���GF��t���i}UQr+����_���{���o��q�(���5\ָ|[�KOpa����q �:�őK�>��\�R�YH�$9�g�w���/J�<��(0{�L��?r����{��i^��[v+.���B�;΄�
7�e�jw��U[A��Ď؈�u�Ϥ�����%��W��P@���Fa�_JX�ݳ�G����؀rG���4���~���s'R�W�2sS������W�D��MaT�I�S�Cğ�oN]�W�Q��(H�I�9�x�3>��AZhVQ��l�w~<{j�S����&�S��NG�d���;7�
�9� ^6�ܴj�W͹[�v���RuZ]׃��=@��"��j���d=��� ��l9-E�1m&י7l�Q���Jh���u��B�4�.p���m�S��$q+���O�W=��K$1@��pA�|�@��M�a~@�OJ�؉���9��	`��(ڲZ�6���
��.+��J��+U	r�4��FU��*�X�����w@z��kՌ7W�ԣ���r�h�d�۸|�x�B����2� ��j�eifr�x���&����=]��h��<9�!��r�9w����ȡp0��OJY R���[�� �̕�G>X�^�ո�c]�}^@��5B6�Q"��5n�<�!�C3��H�w).�~{AO	}�l*�Y���!c��e7��-���]"/���8K�R�����b"�[��-�s4pt*e\s�f��@�w�)(��(W�c�������!��Ц!SRнi0�O�-��E:���T[`�Ls>rB�eI�x��!��:*�U�GHтR�c�#��*����	
-�$z\����ɞ�
��s��B��߄��>��[VK�'���������{C�0V���fqM�A��60��H3J���j���(�QB2L����e�Ω�߼��N�gەMKLr,�R�:Z���l�'Y���?>^�֫��p���W�Xb"�Q?�S����?A�O.�z�h��������&�����r�lB�uG;P�U=�'�+���(/�+?��Dg����� ����������F�p�;���Ww���������KZ�N4G�*��<�xƝ��y/�+r�$��4U�"J�V3��y��ܕ��!aޫ�m��|�,CغLK*���,:'�O��fa�3������m�kɶ!����Ȫx���B�2�B)(�
f��	�l�W�U�E�$�З�]�IL�)w�d�ӽT�6�����Ɓ��)���c:Ro_������/���X@ǐ�{��>B\�14k�h��I�q�kɞ��@V{��f՟����:��v����DD�RL=zU�(b>�t�T���_�/N�^������#�D� eb��o��*h.	�)hke<Қs<�o�;�:+���0���Ơ)�*�P���
��z�U��'ܡ�!I<֫��O|�K�i�	F�:��̵lιmlƱab�6��LbJ����@���o%���X�y��+`�.	+�K�.Cyu]��A�	�3`am|1����� �,Qa�neqM12/.��o������[��M"��D�a�E���p<}��l�7�\���ݟ�^���7z7���[<sV4v��|Y�Z�,j]���;-gs��8�\������x%;L+�h��$#~Uע4f#�6im�:a|o2��Q���5�·���FɊ�ȵ��0w�UW�1��bҎ����\b6.�{k��)#-�"G����(��	Tg���T9���n�E;�cg�1��ʁ����Dr�G��}yv��z���.�|P�Hkj9���~�*U�D9�c�&�/�vr�Sǡ�EB��,cg'�ڇ,��kP�.�Ĭ���.&��ό�[���#��'Ո,#0��޵�m����ˢ��@�H�o9�q{&�]�q�Y��� K���r�b�'��Pj�0�x�����s�nW ��G���j���Bjv�E�`x��z��҈$?�"C|J��jϑX܋$�ا	Թs���  �?��q'z�mt�f����:���X�9����z����"<#�GBG_y�C�l|G?���&>q����*oe����nW|��Z'�n������n�9ɿ'?%�[���Vp�<8Su��7H�h-Mq�4��V&CA*�\^K�K���iЇEC���\��W�3)�Lw�OS`��wvn�+��)�C�z0#l�8���jKV� z�����/���g�ӯ>���&*�駖�B��.I�Z?��5e��@�����r����{������I�Rp�/�S�v����I36�%�2�Z�2�T�uóڡ�@N퐎?E���`n�����Q��3؎"1��{<g�8��j�َc�b��|:��#\�U>vi����$��n�����>&��#�	��H�?:B�pi3�9	���y*�pw�%i��f�f�J��o�Ƿ��`��� ��}7l�w�'1�Y�b����A/2"$Y�?D!q9<��EjXe���6�����N��s�\�挋���k$}x�*+	�6 s�fЍ�1j�1��/r��q�:mw��x�e(�|��y.r��b�PI򡾔r�h��%pA�_�yq�>K��	g1��^���K�p�*�Kճ�.gj���r&?� Y3�ز��e��eΉg������c�)�A���zT|�SslGd ����T)��8�S�Hͪ].��r�IHU ��N�EU���A,�+�2�-t�f ��wv��:}3ZH��u
�E:=�{� �r1���P2��U~��A���aN�b���a�R�f�Y0Y�,&F'}��v��~�/#A�	�~-�Ez�O�x��@qmff�����"�0j������!�v`
�@����+���$�r�:��q�s��5�p����L]���2��e�w%9�Ӹ���ç?��f�t�%h�(~�V��?���
�h<��H|/�~4oHVX��>��&��R-Zt��v���"�����05�aq�G��t������&f�!^w�X�5'06G�^�i&����+�Dr����h�UdgAS��d�.���a��9� ���v? ���渉�ƿ���{W6�΁p�� �7�щ�� ��d3�x��J������{w��誷n�. ��7Q� v���$�]$Y�� ��5�vUXd���Vڿ�}"�D�a{%1����%?�}h��U�#��*"v@�}�����O`'��{�,�{�U�t(�TW������Tm� �o��=�"�IB^h�+�7o�Lr��`*}�T�7�|ĝ7�?�~-�ݪ�Ļ�����s+���q�t���>s|�`Ѡ�� �����כ9�s�B�-j`s��Q6�_h6r�cw-�@B�LP��q7z���
5e���m���0�bkC�����Wzy�84����?�s��g�Q�5�����p洛������'@�J�� x�Pȓ��7�eX�^ʋ�$ډwح��x���I&�M�5-j�鏸}�b����*OÛ=ӑ�]����|�>"��w�\}�#X���u�p��ZdF�u�&�C�W3DE�w+v��>�-Gb�K�`#��@��yQ�G��a��A�)ҋ�!�2أ�j�V�*�'�i���Q�Af�KM�q� �b���h��Mo��& vt�d�-3�ᇨ�y����+��=M�EA̍�C7�bD�}������v����I�Y�f���<}_{5�L�vZ����^��.���P����@j��8�GB�q�����0XKѽ�L�����K�a@��p�)����,�4Az��U�̼/�WW��pC��0ϠD�a^3��ZZ�s�j�(Fm`B��I{8I��_�e	;�e��r�E�f��Õ�j��h;"ܶ�z�g���(���?R1�P��3vK>T�bJ��S�z��J����uGHx&+��H ���5F#�'���1��/��N��F[�`pp��כY��v�Ak$�傍մk6u6Ӷ(���~h��U�8�.�g����%J��E�S��5�0.
a��_BfH�]W{
�e.��"&Vx���Q�&��3ly�pihJ�\����?�x�=�_�?�:{��R&��;���Ht!y�}ƍe2�A��W��4������k2����ط{0=�x��I���Ik��;��ͮ�d1��,��&Yj�Ւ0�o��3�Io��ũW�2�B�gwG}��^�P���ei���v�]:"4�O7�Qo֔w��({콹�<���%1�wR���yz�g��_�Œ5-�\��l��B�/(� �.��Ƣ�L�f�ڊ|�����ƕ��#[uGq�t�ٺ�T��0o�H�h�����Y�#�l�3��C�q��$v>SAup`\��S�D�BW�}�b���{D������$����_��b�����?��W@ǹȹ�N�7���kb2+��0R���]�#�_J<�Bud���h��s*���~�mq�y���';f8�,�sL%��{�w��`B����4�R��Y�ߟ]X݉ۅG����?f]e�jc��V~��ZLo�[��J�@�z��h#z�HE�q������F�f������MQ���#r��+ޙ�!
Q��|檬�M�T�Q�ġv	���e�����!&�������f��*j8�x�_��W����h#�����v*y쀌�3��t�9����4~O��9\d6F�)��42[E��=_?F� ���!�V�U�h�Rbv�-09��x&e("ݩ��廩������~�
\�{��r��=�u�_�|]�÷�>�S⪸�X&������W���x��JZ�:.& �=6h X�Y��s�
�û;G��7������u��-���D��;���������a�j��?��8P/w=���w��Z�1�K^'$���aĸ7���+��&����c$�WY!��O���.z�Q�P#����M�ײ36��+ .�E7�on�S%,b8�1~7������i�Z�w-�b4̘O7Q���~3h+�%&�Abų���ORVmJKќ����}/R�����G3 ��/�p�Yɡ�a��k�O�iLd�g�Ղ�����v/=d~�Pn�7 l��� �T���j�i9�<�� (�A(�pȒ$_J��~����֭���>x�	ݟY�Y���E	԰X�:� ���6��8��������rN��S���2�c�v��@{<�賶L\o�[�&Ydf���4V���e�� sC�������`�+�y�ƌ<�?�`;EP`3�� ��L�B��0��[��'7���;x�=Q��B�!��lB�n��X�>�:���P�K��XZ�98��yہ��m�B�჻V��/g��>������>�e��J8d'"��eQ,rf/x��U�c<0�[��6H��-DU�j[�)�݆$��6I�Z�Z�v�#I�xSgZyMH�?�0��j��w�����7��u>�m#H�E��'���� 6���< �6��dT������f��lcﻅI :�7��X�8$F%K���h�T��I|������k@wx�D0v�Ю@z��ٸ���zI�-j�o#�F�]ө���]%z;�>�L�"�MS��ª����?̳A\�i������y��YS�G �[�3��\桛�SqF�4��c�؏�J"�LԲ�vJ>Q�&���R�P:M�V$�����Su�mވG�xVN���c�I�oʄ<$DL�#m�'��"xK�-����-��Z�*��͎�[����MAxǳt�<��ucW.�M���fs�����պs�_�5#	�	��fƵ�t[M;.x5�<�aA��Ϙ&��� �&����nF�p<�v$I[ݗ�c4O��,�ٸ-e(��7a���w��xI�yZ�{������X�
û�/-ȉ\+��xAH��6���zI�?82.��x��&���3����{{-Pרw2^[������bz^4	�T�d��aP_���<v�NSzڕ�NI�P��k���9t����W��k �*�t-%�����P�%uz��!?�M� �y��-�uY���zY����r&�t����D����Q�*�̾|k�o��D�.��5�#��@0����J(�5&ܟ��vQS+PSͻE�)W���ŷ���!}�gD�b��.���J�&���D[��I��f$EźQ�x�`�W�Ġ|��g�(��R!.�j�MnN��.oHo�GĔ^�<f#�V��7�2���.g:R�P��hzn�J��f�T�L-?c�rI�c.�&w�b���ϣ����=�5Nu��M�9��0���)�)�%�^{���6�f쫊n���U�~�*mpN����^Z2�FA��wjj�O�R�<|%�4�������Ҫ�,�)�~*�TR�v`�68��7m�y���tΑ ����r��~Ѿ@w��d=M��gB�&�S���ΐC��<�ӫ�@i�w)��}�*]�������x�lRQ�����v�i�pZ|b/��	��֪�r8�.���`ɿ2ZvF�NE�e�ެEF��Lli�А�-I0E�
/m�{O ��o��F����W~�5O�A�ǎPl�6d�}Y�N�C+��3,�+�����~�Δ�`�ۻ�[����[#��˥����_{�r�A��w�����J�l6Q�`���
m-�����60(����O�<���y��~Dp�tFs��G����ο&��v$�[�R���2%f�e��QXI�E����Y@��ᾱ;�U��x��$v��#k+]*�u��o�I��H�X�6m��h��i�H� g���U(>T��>�y��{_��Us�f#�~3���4��R ��j"R+TT�5N�N����l[*}[���£�t��B�遵Y���R��C{��-�G�%���b��?��;2k��'�ae�K��#C���
�����x�� �[���vYe\�8-X��>H�͌�!�Ƃ���4��f�S��4G�}`�F�������Q��?�8,��s��PY�F7�����w�a'ߤ0��� 9�X�]�PXA�K��x�X����_驓�t�/ϠoesYS�.]�c�hL�m��X���P�(�#Z#��0йm�5�F���������:'�#�M%d+��vlx��<����0��$�C�g]�n��-YT��<��T萛��c]�q8~?����|�z���/�m�ܼ��tnϼb �gs3�E]���R��`�z�	@:g�۬��{���t#��g��Qko�ęȅŒ�	+���I-���Cg5����Lc]N�+���a��;�Y���\���=e�sBe*ȳ����a����r%5M
ቶ�,-��Qt���w�d��9/�;�D�7�>Y�Od�ځv{yն�P�oU�	�B?[�9@���8�g�8�;ug��wk�5*#��O}���`g�����O��+a��X*
pD�h�'DmdF��!w�@}�/�D�!8���Y����<�J;�F��6�X_��t��p�@���IX��Q޿o�UTeK�n���­C��0�����"��Hۻ(+*�8�vt�3�9qrƊ�d!�Ǿ�}��f�[l���}��BK�8� ������|�-1*�,��92���E=���Ħc��9V�[Wn+У���
I)� ��H��LgH��;� ß�t�y����پ��n5?ӂTI�Rv��'��BA����n30��'b�2`�0��6�%�����W**ql�}9�*��U*�r_�"��Hcөߦh��Ӥ�h��,8y��A�u��u�Q���a<�1�r:�]��O`��\#(��5����P�����@M,D�/����9sy�y|04�cN�S�j��v���:hn�"�]aK %|D��%����ǴaX�jj��5Aγ5���v�p'�9o��a� �m��L@՝��;Yј��;8?�\-�E9�u[�~QşyCpu�$6�� h�G��������9wz�b�L�:d0��n��m/�VV}e.~2��\#�`�N��b�Hh��Q�J��h��i[��//�q ۟�A��R3����8�F��L���H�'�
��@���#�L�u���I(R�D��n��$4��>0�\�YY��U+���F]	�F&zy4��?
�l�.{��u�ڗ�,�A��4�8�m����a����Y��6���~Q�=[jUt��`T��4s���rT��$��;�iRR�JJ����	_�ếHI`B>��K@��T!v$��1�Oç��n8��c�"rT}l�4Z��3Zs����+S�t�\�|#�ۛ_�2��}5�*��MQ�7(Y�i�� �I9���d�+6�Xc�+�7�=ol	��jX��3�|���2��.�"
O��k�~�*�����瑡�U�~�w��ϐ��T����A/�Ǜ� �`� ���g�⪼@�>��"�:&�`��O
��O�R���v�(�d��du/Zͮ'�)�	����CxZ���EYFQQ�6]F>F�V~�CW8?��*eLM}��h��C?$lp11Q�
��H��ز���/|3�6�� y��v"�X��L_��P�.m�Y��������#�'Ǿ�ӧ�t�a2k�x��<p/H���\y,9C;/�<ȯ%�Q�Rp���%�v�BQ�Cl'!	u�Ҕ��ɣ��q�_����QZ�ѷ��0�WX���
06�Wץ�i��fD�g(:�׉F���U)k�"s/��;t'�#��m����h{�xt�K��%-y��O�)��4HέX[�Ӓծ�6Gv	QQ��ZM��b��Ӳo��Ar�P��~�s�tI6�Hvϐ��<y���[u�w�b���Dx��4�m����y��Q�	qq�k�i��J��2~N$_ō��9�пiÔc��i�x����M��h�S�=uӵ:��'$��Mo�ߏ��jcP�� y�F{qs�e������+;�oE�4��*�x�S#��R��AɆY�QLٌ�s��%u6������Ir<X";,|��� ��Iɻ7qg�����Ħ�K�:��ę�x��)̜���@?c�֋[oc�A��F����1a2��D�_ÑCn�eb?}:-SB�G�U&������nU>�^�L�����_�c�S������I��r�C�����fv�ǌN"ģ�D��`RH���^Or���t�Q#�_,�Z�L���a-��J����/���ӗ�Xens�)��r������㚀��jO/-9��3}��²�.�nk[�����`�x�>��lF�
p���ٴ�usGJ�m��к��e�ū�4
`*�j���ҎW~�|�F�ё*'z�"p<��ʜ 8fw�,�{�N3��L�1E����d|:*��QpnRޡ0�� jT�%����	9�j��p�!\���^Uj��p�I�$��$q"c�ۡ��,�?�9@�@�A聗���9��
�6"��
����d-��h�o��{eY3˝݃�3*��,��%�>�˚����ÿ����%��	.�5�yS��bq2�x�ǹ�۞k�X4PJ]��P����Z�^d�P�r��[4��&��"�=®�����B�h3��e�m=��:˓}?FC\�f����,���C���`U���ڌ�2� �p��"1�,�Uk����*�p�+H��,�a�R	̣�
�B�@��$��~b��������b����ͺBK��f��G[C1�Y�}�3��������;�0���D���#�n�1����&���m��X��4"`:n�1&�Y��_����/�2�.u��������?�ntհu�p���i�Zq����{W��f�x��.̳S���B�#��#걾bP��EgP�Ԙ[0� �q���կ�����m��kD�!Q�鋙垪P��͠�Qz�(P��}�?0�5bG<�`A�G�N2��SF�e��O7�� �p����1ʪ�]W�p;C*�]�h����L�Z/t��	���"	?�1fO_Ț���U 	=�Pa�.	����D�����&�8���V.|�kщ�q��\_a�Ω��N
�4#��[C�$W����J�O&�:�+	-�OZ�k�nDQnW5�xF��S/�.����q#l������c��o�o,�y���[$
H�>�F�^k�1�����ٛQ}������A�^j]m���܀@�cN��,jr��Ϝƨ=/T��x�zp���2��*!Z��o�voO�9ri۪oV��-�����oJ?cS�"��ʿ���Y��I��t��"�a�f1��\�x����ďK2ve.�D��*sߙ>��$u�x�|�c�fJe����+)�gN�^I=PH�sK�wх�?H���,V��;�1צՕ�2�`�\��	�\^�n���1�\����v�8���k��1���1Q�O�,����!�6HΨ@��c�n���	X*�ސ���nSz��;��W�F3� !���J��^\�nU�4H�yp�|{k=/�x����S	����d�ު꓄~���tĶt�Phs�J	�rv�q�lFT �֨���]�K_��v�Yi��q`�gcX�%<��TW�ֆ�&���������3d�{R�pM�|�cn��ɸ�?���r�OI�b��J7cڍ�%y��������X����{��1���j�)�-�B�L}c��K�5��9��*7nE���=P�L[�q�
���O�~ۥ"
&"���ꕊ[�]���X�s�:ϋ�g��AD��D(����(�c 	�)�u�S����h�R�W#��$�%nѲ4�%*#�����<$&k`��!$�fq�y�ܷ�iȟ~po�=Dq
�A�Mzn���@II�i�~���;�m�	�&A�>k�Jx:<��_�{�'6�
R�+�`^xU3:9g�g�	mMa)q�(�s�][@�
:fցT�2�Y[������ߪ�:�� �D.��=Y@(-��v���Qr'��t��%�¦JORe�����l+�5U,���"a L_N���X"�O�X�NC�]e~�9�x#]]҃�Mx��C��j�zs��h������u���r��.)�]�i����Wl�z��/�ك\�H�F�73"^�M�aV������i��u!-Id]�x�>y�� ����c1�@��DLӔ҂E�0�֤�ћ�ypviێ�����!�	��h��t�y�*�~�f(��6GzU�_m���P}RQ��^ߒ=$I�n��-\�D��C����G�Z����Йbh�
.8��4�����/`�m�E�GOp���:��9���D�k�Q��>&0��q���朝H��*�����d��N��8V��� 鈛m|.�1M��8;�U+�[�������c���t6.��pE��q�@%��g'4ɲ���
P>�%�$���I�� Ǳb<��]���	zL�C��̱�S"��P���ɯ׹��*�J��wp3
լ��F�$�a�&���gi
(�[B
Ɋ;l׊�x�on�:�t_L#B�9h���R�{)��>G��Ǵ{4`�ֆ!��B<�g���>���1Ie1SX���>_]�[W#�J��(�����������q8��Xd��@��X=�+ܫq�kX9����-j�:aW��E!�K
P��)]?5�`7�p*�ڙdhx�0�gu�PN��f��FH���B��%���<��x.XMtt-'��^��E���zŸ2A�ws[hD�MC�9�>�M6bD���լaS�����p�Y�����y��M��o��eu�C�eG���ۂ8)�5[������ƒ��HbP�Tm<<Ϟ�e�s<�2�-��'�zȜk{��<L��r��QbU����掾��;���l��bq��Xb��猭������Z��#�q����nM�-Σ�i���d��*u-P,�ά�@X�xi{�[�g�+�+��6>�΁��ϥq�(<�vf�q������A�I���I���q)��_/�WMe݁6P�G�W�a�J��6���� h�BW�s��I#l�ߵ��{b�Ώ,|�c�ؙ��Y��B�$$��)��+�&_����^gbX��
�����a�y�2!�rp���d]�"�	j}���*b��pN 0
��u�Cu��[���Ww�	(�W�A .{7���`=�d���1��&�{�7'�mZ�qfN�P1v���]�^�?a�0H ED��L=o�+H,��Ė+;���s���BdȝJ��SV{aHo4�Ĩ�-�#����o~��~����H�>H�_���#����H�&ԟႩ�m��~]����񚈗�� 8��g(%ĕ������wS�A��-6�WFC��u�yV�#��'�O��t
i�����{��3�7��B�%�duv�lL�/���(�uh-N��c�����ŀ��!��=�L� �׃���jh�I�rҎ52g��F(�v��h~��ع�i_xB�4!�B���n�^O}dY�Ae2�����./�B3E�:$��/�-�(aN���B@5���}Ouw��Ķ�H0�)��s�oF�j�0">܌ߚA��3�eA��<>;F,G�2��;�-�?��6��o����It-�a+=_x�:`�C3Z�*~ƫ;��My��K��Up��R�;���^��C����$��x#�T4��P�keQ}��n����nŇ7@
����q�,ف"2����1��B������钓���#��T�N8~w8�lԅ�ż�'�ќX��)UՊ秬tA�t�cH��Bׁ�xu�Y��|_������Ը �̲(��$��m�c$���v�*��}��.��@��~����2��A���X��/tUg��3,���'7�����k����0�F�M��#�&QĐ4F�[�F']�k���ڿ�tn�k���&�Cz��e�������]��q�A�#����ǲC:���a���r��z������Ő3ʛYh�CԹƏ�����2��{�h&��r�����σ�U�.2?ؖs�4�AI�r<���7�|�"8�qn+�8E�{�Sꠊ�nr�./^~F������ذ{��OE:�����^PΈP��j9��ڠ�W�h*��TVjI(�"�ڵ2Oo����f=��N��V ,*	՝u��]NT�ell-p���^�^�`�cn;�[�cz`C|���o���+�O]�n�?H�7Sp�ܟɰ�<b��f��HȺ1b ��J:�7HSٕ�r_�хv�$ȁ�t�]Ͱv(�8����B����
WKh�x�uc^��������~���6"M�]}�mm������t��	�7��f�Z�s�|�x*��7�����֛X���]B)[��F}�!i�c���]PZeM�&e8V�[' ~a��0��˲.*�lŹ	���c�EکZg�E�7���*��1׵�̰{g�H�1�<�x��Nn�K�`^�� j�)#&o�� ]�Uv��X57ćQᬸ���\�͏��-�Ip�Vg��P��ns���r���↲6ٛ�� ��u�'����B^����W$$����?k8b�v=V�V)�/��&iW�R\�����k{y_�}[�/���u00���3& ��X�#-U>5]�~� d_q�a^���wV�L��:�7��jTW����g@8(v���<��VF9�ذ�c]Sf�f���^X.���1���'桁�7.4���!��6]9��*k�)7w{8"�6~5�V1\� ����%�����Q_�<�:�m��V^�{`�Vϳkd�'�m$\�����������.�t;/�¤Cg��$!}�P�3@�ȕl/��\ZE8�Q�m�)���\źO�U�e��ԉ;Y�y[�㪳��}���ژ?9b�J�e�kY.eE�"�2���^"]��;��س�:%v������l@r'ICD��0�����& ��苷���y96��?�t��V��_���T$��G�7_F�[_���<��ȉ��NTg�h��f(�5M(�8s��G�����<�a�,J0jI�����Ɋ��K��m�D�k16n�-�-bb���7�)_B"lI��صqI����AV��*`�[�b��-R.)�uf��Bh�cݯ����oM^a��c��y��(v�֧	-}�wQ ��@����C�i����S���.���=�0��̼
{�j`]IA>��Ue7/
�)Y��%����4�?��j��z"O5z>6h�F"~4�l�5-�,�-d��=X�k���HU�j�@24�2�(��ƞ�n�i'�y�B����C�����
B��$����rdQ�QA��(�tcx��S�4S�n�@���������'�`��͖�j����ٶ��=�����5�<�Id����aF4M؆�',7�\y�m����{��\+�)����(�!>�Y�g�0�-�N��ٟ�ő�������������ޗ��+�M�o1�� >�p+>�Ii�sQ6zq��g�eB�̔��p��wu}���|��b�k$o���n�|���4���8�zE��4��MM���u�Q2҉��i�&���$]�xW�C?��:-<mK�=#�o���W�!�<�J��鳘�Fb /˾��0��v@.�CR�鲸,�����r�%��9�2�:����#!��=J#�c�wi�&���!�$�����U\�8�>la{Z�W���$�;���D�]��0o���w?��)�$�GT���6�_|�.[��kTz<��Q�`O�]�o�����:,%.%����)�����k!��=��ı{��#�HY×X'[f�{��Jޘ�Ɲ�ą%����'l�T7p���Z���0�|%Ɖ�lR�T�.�EFh�~(ye�i�MwIO�7���=��+�3� �B�_��ѯ\=@�C�4m�{�B���R��;G���[C�1����_�Ct����W��E�pU�Q�EVFT8'"�����$o&M�L���ymµ�L�9��K�OD��"���Q���]ٚ���F�#�j,�dR��]bW�(�I���'4�DOX����J�0  ��|����S_C4'0#Z��q�ʑ9_���Y�!V��:���H6��-2J���~Q�#-����-0��?����(>��a��YF��#�&`�3E��w�թx/���z<�+.2���*��j/�{	}�t���X3sK&(�s����!���Q�b��G���C:$�׫Y��wyu��y�v��*�����Z^!�{��%��@DyT�l�k�9�y�B��6�;(/&��Ã�{%=� \��!$�߆��0���=��m�y����<z�B�"���R!Ȋd|7Q" �$ш�f�;��y�A�qI�[�ϵO֐��gp���
w�n��0"�#���4���+与-Qcm%����k4�t'�`�Ӫl����;��lG���+�ޘ�"~��͑`��B�`?��o��.��u�V�x�_Z%�	X�� 5y�N�5�@p�*Q�7�\Նv�&З}�Feu����B�2�a���5>z,@@M�؁gv5�ںJ�d��"݆Ҩc��yOߺ��Ct�����E���a堞�a Y������
elx���!;񀸈N��$�<��r༉��-�рV��2�w�H�� =�Ƚ�l�'շEl���~`1N�G�N��̀�G�l��u�Ƃ���!�^�{3aM���q�WXM��c�����5X�7U�z��?I�G�%岱�����N������u�U�C5a1C�L�h̑	8�!���4�)�
��4��3[��Jr�D;���{ŭ�YFk���ǳ�s�d9Q���`�A���Qœ� 𔠴A��f�H�Y@���6U�p%P|.��Yv�\F�e>jI��Q���`��=6g�Q9��(�ߖһX�_~�.�Б�t11�.w�ֳV��È8 N�����=�;T~'%�o銍���l1�Zb�xM����!R�k����ͬ�l��)иd2���Ĝc%l��hWm��aa�Ŵ�����4;�rbt��ߘ2pwt�D�-��b�#@Z����v̔�H ���I�[My��VA�c) %GN3�q<���ŇR!���qD5��0r����F["�@;�8hy�p^�e.��;i������#�y툡���fϴ��6��)�_�k{�@p��s&�`C�-\S���#��C���u���"���Z&���jB�h@��=��ǅ��H� �2���H�}�h�M��M8�'L�'d����:���<�Ɨ����_�Q�5�4VM����E1�E"�јON+9� � �#v_e
,��w��'Ԇ�hz����ί%�!���������ZA�P��՘N��߃��JhJ�Ď�(���`�TuV~ir+��
YzD��ο����`�v>�s�l��\�n�� �n�$�������SDL��N�T�Ƌ�S�*����nR�M�}�࠺>.{�q=H!�4 WP�����g<B$��O	�ԛ�΀ޤc�"��o��wТ�p|�Ґ:��/-a��`b�`7��ui�U�$?������Sܰ�V/���B�.�N�J�`���L��:.$=���/=TIS��	��oI|l(U"�K�	U�߭����7W��O�VJ �|�!۴gr�[�5⫻.'���\"��t2/�(�=����Y���A"`>����8pմ��ݫ7kX*NL~Ƣ�����?(5Kd ,Ά�x�$rB�s��r ��_�c�O~oi�Ld.��b!^�!�K�]��{�̈́��v��>,5���Uw���4l�����ur,r��^#��P4/}d��#A�"+��T��9�Ij�����\I�'L���=��`�r�Oos����6O���-4�#B�߹`w���W=�@yn�$'����m'�2l�䐮(b!�}��<�4j�^׉��c�����!-�!��N������|u��
a����_N8�E��G�DR95z���Nܮ�T��������E/�"���Z܊�	
��o�I)E�]K/r|�=� 8㦊�{��
�V�
7��@`����.�S)�R6]b�Cs���|O��NE�/��7�6��nz��/�:�P�����p�Q���;�Z����>��8�Ӕ���}��.����l.K�c�}�͕��lUa KL�ݥ�J�K/�k<>����j�>�t">n
��Z�,:;=������c���7L�:�⓾Y}TN�n«��"�X�i^ ����X ����=NTr��7���j(�yRޣ ��g���OK���?`�����A}?6�<�������x.Y�Z�<j~ UF��(c6���6��a���L���T�k����(��i?Sh�Tod�p����Mo�Ѳ��i%��Rw��:J4 P�G�i�LE��R�G��>N�j�DI��IQ��<�VK�q%���ȧй�S�	A�Ao�ʌԗo�r�X1�M�Ɗ���5;��Q2ݝ(6XU:oR\L�w����}%�d~ޅ���Gc��	��W6g�-�Y=NN�]��Z�h��6A1�մ�JY-����jG{�G������_2c� c�E��=�I6�c�fCh�P���7�̰����VcI}�]�3|Dx%�?�C/�2=�pFTc�R/�-��t?ڪ�&�k��L���$��w�`y��޴�6T�����)��V<�~#��p*�Q����]QC���M�
��l��@%���x�����Ot�d��0o��n<���>���V)�]Qe8�c�α�h	o�V��肊��{�}*�x4 T��e8lT�!MN4=�s���;tfK쳻���\]�]ftZ�H�̨a6&=��٘��n�����3��5* ������kz����%c�
`fPF�S]ԥy��d78"���.��<�Fq�ևH"���ʪ�B�a]a���.��JQh:;>.�;��@��b!�/�r�PJ�C�XCC��2�9�5ʹۆ�RE��lo�!ġ�Px�_�/�W��Q7�bQq���)v1����%����I���dylr��l`
VU�pO�7ty~I:��o�Uu^+^�j���8�aR�Q˛��v�P3 ʟA�\��>m��V��j�$��r����x63�X*(	3� ����22�f��d"�T�� g70oXV�qp|hZ4b�"�T��� ���-�r����,�L���FEm��85��ٌ`�-��O�$#v�����q[Z�9��kT�A�MT��gI\CP���"�!�����nRq�{fǄ��R��B���q>3r���6�4��q�<|~ �S�m�_�1n��jf238`�ɩ ��թ�#�%e��p����f�9Pr����^ڪ^yP����]�p�ȀD��s�Óf���[:+�iZ�C��Հ��x�8�����_�-aB^�.Y�$=����u['�����^aT�2w_�Ef�O�xt���������fZ1yc��F��=)��"�4$c:�G'ZN�������t�e�����k���%��:��-���r%��ŭ�Z.S��d���\�kt��@�Ō����$�Q�W"r���$�p�VL-���:�2����gGI�Km�����a��H�*L�b��pk������gͬ=���U���4*��xP:�\��1�W��wz�D��|±N���%��.��Mw�\&M��*�*�f�.ֺN��b�9���A��;���s�{�ؼ��_�I:���1B'��*�� #��|zMH����[���{L�9��-�}�s��|��c���o��o�E��췛���= ����t�!��������Cb���O#M<'����93�t�촱Y$8����}<kI��1Ui�|S×H�)-�sּ>`T
�ިJ]�ۙzYJ�Y�-�<��@R.���58x�tVA�
Uƞ!��p�4�1�����8k�6���r~j�����xgA���4�Ԙ�Ԍ�_��F�t���>��jf
x)\V��>V��F� ���rS�w5��A4����d����]������f�|vR�T�L�dm� �p�7{>�/�Y���[�������>p*�+s�N�]��H�������r��qNĹ1!��~$Q����:��9�2��0�LשO1�����Wuc"C�&�O�Y��J�pINp�=\��у�o��B>E]�&~وI+���:��{7P���Z�\��bJ#x���<�xaA�K�z��bc�1��Bp��c�y�0����;�,�_����W�ێ7���VPN&x�I�� σ%=f�Y\����f�j)
G�YBAFLm���� ��N�%v��Oy�N �5��;��薈%B�$����f4�z�uxu��z&����t�0#U���
��2q�6&������?��rt`Yk=����F��ZO�S�i�X;W�J�r�JuE$��G��F�=�s���^J�q)n�;v�>"�$''�O��#���7\�7���Z��5���������d���}8n 퉳�Y#b��)1��.��3E�kT]�~m��0�贇4#���
L��z��f�r�C�I��i�a��,�R^epTP��Za�=ߡId��� 혠���:�} "�7��(��9�/���C=�uƀb�Q�6�&@'����;�3��6;=>� ���y}U6�3��GFs�zɵ��`�>A�t�7�|����)��CER�ǖ�a��ٯĿ�z�OIrKk��V"y���ԛ����ɺ܊����0n5ѧNc��D��ZH�ɨ{Vw+�7;��=~�����|D�"�~E˕O����W>����>���r��+nֲqؾDd��$Y=H�'?8�� )Bk�2@7)(	��ʝS ��X��Aޠie0�k=��dy;?7���g�F7kJ��$�}'���r�������Nix�%2H)�B�6���M�L��a�7^�:����ir@>y[��̆��{��h˓�B�Xw��L�
�0FI�a�%����(�]��$��rH)�tC`��Z������u� d��E�iB��o��:ޢrȑ�)垈#�H���B�[�8Bi�1��U�-���~G#I�*�lh���4J��	x�2/�a���;�Zx9�	_����L��r��O#P����:��t��u���i��.�L�(^�7�@D�T���xN�!ʰ�ڟI����׾�9|qſ��&i޿�2����!.cO���NU(����AhF�n��m� �pݒ#���������'���\�����w,?��g2����L��%�0���b�f��&&ZY�1�z��vR�ڬ&��S�P�H�6�3g���?e��ϋ��a�S|��S�2�v��+�J��jT1�J�Lc-D�(b�=�@�!3�%j
�T�	�C%S����Y�.jʡ��}������ϟR��{{�u���s}���_���]'"̸��	)�t[������Ru'�kMd�ˆx�>B1���d�s����0	*"�`�K�..F�%Z �@�v1NA�=Sg�{����t/�@;G�6�N��jͺ~Ͻ�.����cF��H��#6+���^H��f��̷|4�G�Qo&�'�v���ȼ�ps�I�J�^�t�i��5&d�H� F���>!֨L��ļ)�I�;GĹ�A�t;��Tj�9���/H�#L������<��}��,�8���Űۑ�*o0�*��;���N)�N�T uI�c�M���E�b��E;zI<5o����|qƤo�� ���p�`�π���צ7�+�@�0j>�b��dCO��8~\؎���r7����d>^�Y�c�:�G2�oOm{@��Y?�da���H���Z�m,�] l$?qG�]����Jx��� E�ߴe����
	�&~�u����u�=�����$��d��GŅI�T(o�ɉ��8E�G���j�y豀W�}"��mR�)�Ԭ�Vu)�}h��[���{,fԧ��D�ݓ"��j8e"��g�W��c:{s��V\��/���b�K�,^���ݪ���hT�o߈)ϰ��W�����NQ�+��I~�h���4O�w�y��7��Z�w
�;� �̞^X�-���*��űS��%S#�|_�ñ^ a�U
2il
��	��孵ѓ�>���֟{����L�Љ�%;͛�HhI��T�]�42�_���)!IU�<&R�W�0o���0�Dtl���6��՗x�#��5{�p����m�E��σ���*8.wwJ5^N�?i�WF�oW<�(H��Ij�.���C%�+g�#�A��G�����Թ�&O5��*�$/$T����,]%�.z��E�fX+����3M! ��z7s��w�^-/�7ݏj�xlQ�;:q�[a`a�n�KnD��=!cb`xS���Ա����(2�`����ޟA�\(�O�T �c�;�}?�3K��13��m��/�;y	f�خ��)�m��T7� L����e��i���W/}��� �Q`^��N^�����삨��~�� �h_#���zD���?��L}��ޅ�(�+9��ii��)*.�.%EV�&>��I������ Y0������5�'_�L�u`���;[$~{/R �'/��' 	2}⦪/��t�%K�!ؚb+��B�<ƻ��W����H�$��x��0�Dy��k��I���G<{�$0^���[���δm�D;OpPZ0�^����uRV�]�e��Q�j��P2�br�@2�3��%�<5��O��^�{+e�v $�X��+��&��S
Ny6ν+�*z^?��hܦO����e��	�<7�**�ʒA ܦ�ӒU\����֮�)}v����藡�f���4l�/�4����'&�d�.�.�����x�{�o�Q0&�P�Ip��������8�7<�>Ig�i� B�]A���g�o_K��'.!_��%�h�>b�ۭ�Y oy�J�c�,�%�|I���G�g�́OPD��W����1P�4�6H��������呤��cY`|T�� 0�n��v�p�dB��|;���ʔz��.䩌���1X`������h���3,�, r�Vv�<�����9�K�}��[��k�!��W���~�I�� ��Uޅ��O8���@�r������;x}n ����<PF�?JDL�Uj7%�/H�x�t�Fh5���&����֊N�2拻��p�?��* >7��bs�-Y�Pb�2T�֔�vҒ�A5M��+j�x�M��`�	Ś�u�!G���	�V�k*��3���i��e�p_!������{_VA<&MBϖ�e�C�U���������riޒ�M�<w�L	D���Q���Y%0���+���V�~��� {�fԫ������"���/l�/����K}ʈ���L���:��K���n@���ߟ��v��R̕;Lt�I��sEf��xf���
w�i����v�V��nG���2�r5	��)"���T[j}��`�k/<c�[�Pn6�1��9��ރ2r%�$�tb�B�����-�^1haQ+U��Y"a � ��rĖ��Us$$�W��g����p�]a��n�j�>�S�e�X��.��k���۱?OKC�6�FW��.�RK*5�W����3��zS�/�'�l�1ݐ�	]�������%0���ǵ���Ν�.��j����:���>��M�5�X;tD���@2�����o]qn5�+�9Nߔ��?<倿�r"J�^ٙ��ܡ�T��������Z	��a�AC��z� A��>y�U�^�#7��}[q�p^�=Y��
<�y{��y["0*����n����b�!� >_`p�q�	Rڬr)�[�l$S,��2�t�q)i��Z��8��xcr�F&�i]c�͗�=�rJ�4���v:���D�7��}YJ��v�'���'s,*ӨL��`�6v`���H}�$ę��}�F���q|n�_7�x)�)> ���`j�m_u�<\��9�ˊh��#p�ۖ
��z�x��K��W%k��,'��R�\��`_Yб����~���+�~��.%B8�7ؑ�P�(�x/%'Lơ>)b\�gn��	v��0��b���O{"O���p����r�ӄsqA��ۚ9����d�&+��VX�Z��{e��9����A�Z����>��<��S�+ڬ&�$�\�37�hg_xu;�ش�������b�ӗȣǌ�]K���	3�y>��9;~^q0�	V�v`/a��<�:-Y7�ssݳ���E4Y�h�0�f�#�/:�\g�S���@@�0�����մ�@s�����^��G��m������ς<J�c�ӄ?kr<[���K�:?����P�3����G*�PbKcW��4Jo!�#�e�n�I�ȵ$��+t.7]%�%��q�kq�A�:k`�����I�8RH�5��lf��&F� c_�|_�_C�ךS;�o���|�����1庪�iɡ�`��uE�J�C�e!+ӌI,>��|��EA'	p�|e�ޓ3�lD�f5"��W �Ͻ%�aPm�m잛��*�6��*7���l��Ə�mS�`�܁��L5������bS��Я*i��g�9}�] b���Ƌև���w�A��UE
�Sn��i�����8f�KQKh"��TE��Y(�y���Y�T�v�� _����czO�"��U�u�XV�G��}Y'�K��S�ɍCO�v&��� 5��]���l6�^��	�����#�Y�b̏�A�y�8A��|�Q�A���'2L��#��� A(n@�A�v�8(�|�j����
	�gY�%~fj����I�����	�nq��Ь�,�d�M�fC��w3��M�C존�ܤ�<b���6;R�޵T��%ivjp��գ⸭$��nܓyPb��p��u�D�_�4�����_ѝ�f��;,�U,®����(��KԷ��z�ρ�'��r��P�v��+%o�TL�{�#�����%�ESHy��b6��ѫy$����ϣK̐�s���
ERq�e�4^u�ɜ�mFŊX���Ibŋ�����\�Z�ֆEĀ�9-�`h��Q���`r���p]Y&��4k?�\�xҬ�9j����Z�����t��Ҙ
��G� V������Ti ,6��|��Č��Y��J+��8����yGm��gn��Q��>�l&ʩQs}�,7vZ��������A�ٻ0͡�ZP^��]���R~M;-z��n�^�ƏQ�`��5�w/��������� 09�і�-:��O��D[�_!к7؂��Q�Y2�
��YW�������'�hEh��I�́�$oK����y���-&��*��v{L�:I:�O���L�%�S*9&6�_k�t�-I-=-Lf�-V�F5h{/���� �v)g�7w��WF�cG0�����ɴ?(Y��9̏\E�i�\O�D$ۄ��ߣ�{t=E����$�^���hk�r,��P9����]v�� �#�	>���μg���S��'П�Uβuk��~|�~:�颮�*�/�~ɒS�IR$d��l���Q�rt� �f�7��a%�Չ�|MP�ԝg��q���p�	NE���J�T��H�e;����@_U�L��}z򤡚i��~SzU�es2��ُt� ",y��`�i�ʻK[׃��a@�+z�����H!��(��e`.���z�޶%)Ya�;l�����~�njf��k ��>��i�'ڪ�DLoN,3&��j~O_�}�~dYo�=�7��t��ʨw�:B��2�����U�_2l����*�9���vz(�G|�!T������� �9�8�����G���4��5���(�v��U���I���-j�y��D�9rq�YX-c�h9��vm�~ŐB�c����-!c ~5a����:��`���!c	T'c��F<���di{���Ay��Ƚ(�0�ˣd�e���nܼu������pk)Z��.dx�:t[��ݳ�K��B�awr�_s�:c�s!�-�]I�nG���g�z]�\v��(uEEhR�sd�"�M�.n(y��']��EZ���[=��Z��"�%�N]ਜ���T�,&ڷe0k,~�1�H�XcE�Hγ��r4��c�A	�W�W�l3p�g ��=׻��)d�]����Rm80����>:E��o��T/
ѶC\��|���7�NE?tD�^!�������9���7�4j�F$��C*���#qg]����+�?:��+O;es9�u҂���PÑ*P��PC�p��� "�rɈze5W�m�pC�(�-�tz#EO�xba�'>%�������Ӗ��wEN�_��݃�D �R�$�̟>����5ĥ ��77=&�ӏ��	N�-�k��:(mI��"9��VP��T�<�Wo�,�b��A���k���P�ت��\�3��g�Q&���t3���^͢R�AF9�ew)[e��).�p������Y��D��!J9g�Y'�,���#"�?q�P `>��*���و���b��O)YYe��b�I����
�A*��3�U9�R"�O� ���L�xַy�X1�z=�AU��0X�������_V�l�t70�_��,þD�Ϗ�-b6Gd���.��%}@���Cb�y�7��Ms<u�ͣ�t�r��N\;�<���!{
�K9��d"��F9��<J��v�$���i�q�|AZ��v���9`��Z�+�X��%d&��etR�o_c�1����S�48��_`m�L�Y�
�9�n w3an������e�:QtRmи)���gw�T�qJ��G{�w�* �Td)�~�mRY�b����g-ƀ&�{sWqxwoC�3�S�/���hR/{.�" ���l��e�y��ֿ��s���+��T�2��)��ׄ�&��q�"*ALF���^�{���&B�"W�DD�;��R��4���EyT� �ߟ\9��+=gy��c밄�!������b�-�w�����=S���2ɛ��#��T#�)p��L$�D�Mnwi��;��=��>�K��zq�)����EHVe�`���kB����w��P����9I�V	�3Sc���3�|�W�d6�����5������\��Ƞ�}_A�P$Q����5��:���v/=��>	˙I��h��k���� ����}�!��PL�Q]$W�	#���cBl�PN�%>�א���3���*�
$�mt�����T��t���
���z�d��_s���i�O��'.��.B(�m�-�2�eb]�7;kr�xJܸ�%]1d%#�	H�U~bv�s~[O�۩����|(�J� �8�x��'�#�]d�WM��=�,���"�K��h����ȗk5��}���"�'g�8����4��4��~o M�)I����?m���Xq�3!�ڒ�� ߛ`�]b����n���Cx�0/F�}���A}o(hPŅ��"`�*Fy��n���X��L���}X�v�X���9�m��N?�V�� s�{�z��b�1�����`2����c��/��T��B6�
"2kZT�3��%����oBwn��`�]�5=6����`�i�☆H�(�>l�|�N�e�S+������}�>�e�}�%βWp�K9,�	8]��u7���A�i�>���It�*%�!��T$|�"\���:�C� �7��:�z�����!mM5�$N<ސ�Da�.�i<;�����74f���c�!Q�MG�D��ɬ��b���P}��dKz���߁/���O�X�b#`���%��-�H��)�,C��`�A�~*�6as͂�[�$Ns���I�M�������e V�f|>�MuݚA�n8�vTA���x��wMR��FJ
%�b��!!է�Oß����G{�����G�-�1,64��a�S�����g��F#�I�,�'m�/�_ț��>�"�ڗ����v!O,�	����9�=��<����{�QG_D�G�k�	�t�����>`&����}��Ti[��C�P^S
�z�Ҳh��O`͍�x��F>�.X�x[��{���B�ڸB;>�>��&�p$�`�����\�@�(��y����+�Ŕ+�6�H�7���f�POd��#�����|��mGԉ������E�{>������1�
P�H��P��TOݛ��/\دj��wO-	��d��~9nl*[6S�M(�l�K�sk�	�wJ��*s�=YL�6� ���b���s��Eff��lF�����?vNZ�q���I�b(�$>�B6O&��� �/�`��z�oMX���.[�^{Z�4�rZ�r�2�QtH�f�-��C�^]շ4��}e�|I�M�n�`�Izhilq7�N�W{Su���}b#ȇ���߈U�GR�<`�t��@к�Q&|R _ܸ_%�2ЋO-�mJ�0��b�n$ط��KD�����qX~���5�3U�~t��8�kvt�b�`m�6J��2����	�0Ǽ��l)�jq��G�'�����d��i��K�5�_B�?�Ϲ���X�!����*
Oܼ#���g�V�V-��Lg	�]�܌dy�)k��=���.V|����&ch�w��yά�Wq�v���a �I��^��`���[�F��Ռ��:$���?�jx�+9F솛r�tr *����%J�'"N���W�!�}�f1a2�5�L�+:�/��Z�C��<�#z ��鱫D$.�z����0OF-�V̤{��Ų\=ig����aY�޿K��q�lV��qDZݯ��zg>��&5Z�	d0�Ϯ��&vZ64�0?�ܚ��6-p3ӕ�@�O�i�5Vϰ�3���ɽ�iv����x�ڂq�h� �߸@��������<ˉӠ�Y����Gu\�W |�qHb�2P��cE����[jj�˜�1t�/�59��V|�2�d����c�r��*�m�Է�<w{h����K�m2%�>?@P���W5utQ��P�m�qY��T�"RL ��`�l������5�b^��{U���?y��;8(��{�"�uB���$S���X��a�_����	h�����qAb����$�KJ�	�_3�,�|��]��5Ȋz�3�3;�x�m�؏�!���}�������; �1o>tb��O�4mIڬ�L�9iɲ/�0�ٓ����I��s`-m�Q�02G-���0 �M����땤�:f �p�B�� �� Bzy�"C��~E��_Zfc-`�b�(�Xߑ�� bn�D��S��b�QZ;ej�ݷ��Z����b뱝^ȧyxٸ�5I,F�֣p��p����ʶ��+{�%\[Ġ�{2J����3P�J�����Axɩ	��Q�y�ݤ��ŮtB�u�ǎ��$=@����~u�k����,�x9�?��,M�
K��]�Ðl�����9f��E�
�-����T�a�n��\��w�V��>�\gu�)Ȝ�ΩU-��U<VL�h�>�ׄwfC�i�E�W#�<ޮzs�;Oڝ����K�5�*�㜚8���@��A�ǆ�<�G���Ù�e��>>J� ;\m�H��g �퟾aE������@��"�����4�\�Uq�V�����~�]�Ea�n�t��:�{ Wd
M�?����?��Ndt��R|=�a6A��M�1�-�$�ׁ�lj0�F8=d�:��U]5�se���oi��t����(��ً��xe,B�����6ެ^��6�G��5b(-I���&G?���J�1��|�<����a��ԥ�z�P��E�t��I���kͩ+���Us�q��Kˍ0���'�8�~��a;�+�=H����x�S
S�Q����:y��	'&X��lFS�w��1E�E��[?nR�_�xJaߡl��Dt�J$_.���qf�0�]�y����Mx�fޣM`�_᙮{�vN[Wv��sm�͊e����;H �\\'��Rp��j7�0���M������|������,=K�w��Io���ն�o�e��%N�4�rui<�ȴ�>��ЖF*���̇ �熢4�N��	AR.�ս�>f���:���,f��{6��1�Eà�Q�a��=�5߃L, �9�k���Ru7�	�?%0g�dZNj��8\Fǳ
Ѝ��9"J:����\�gJ��2�8�p(~;��^3�:4�(	���Z(EU])���B{��������؉u\AH��Li�6��7������b���A�0����'�x�+N�{�`Id*��0�O��Y��H"%<��p*�e_�1{�+o����tAםx �Zc#���*Z:��$đf`-��Qܒ]�^(xS�6�{���L�IN��>e�9��3)f��x���<j���'�Fw�C��QJ�(Mٍ Z��eVbr&�����,�$v7��V��cɳJ��^��]���]2��G~��=i��ъ�(��>�ujU�A���LEz��]�c U-��*���V	�f���x�\ ������h��+��7a�J�E�����z��R� �g}ߐ<X����u �>ڪ�Q�F��WF�^��a�[Ѐ|(�p�>��樢ģ�j#tE$�Rʯ^�QZq�^ܑ��_��+���VC5�;�(.7�g)%�d	46��wV�V[/r;���nfb��+DS�ǝ�h��<v��*��)�`��4�B�(?a���Y�B�O4m��� ��T�5�� �����ZS}�"ȩD����Uu�5�z

�َ�*vO`6�^�8N� KJ�<������ޮ���򻦵��x�9m�TI#�x�v�ӏv�xPA�`��o58���:��ц�t����ܺ~�3�g�s�?m�!XbI7�+�&�����pdl���g�2��l9�?���4�8�`��(ﱝ�X��y�/iF� sY�5�.j=�����o���=������ֆ0��u�#�J��2mu�Y�����t�O�5�k�j*Qg�g�n�C,��2$,[0�DU7�0��,2!���ϫf�՘��Sې�mt�i���b���d]����7����*R��n^���c�L����+���:2��j�2�V�Y2�7d��R�c˅3�<�x׵ ��¬����t�r�9E�X"�	dnI�0g�LV��	�C�!w-f�	��܏c�x���,�9���7�tm�ۺ<n��@<2�W�yU��i�č���[��H��ڭ���HID�Y\��&���IU[<�x�9�@�.0��if���);;ϡ��د7�{������yma�@�8b�%ಾ{y���bP߱C�l���\�iWjfQM���̥^���0�O�_�8��^���%��Q�Ċއz5�U���P��}k�F~��A?�6�`�(���T-um[��T�)���'�<rHkFV2jz��"��E�R�ݨͩ���W��N���B��]G���`��2��jւ��^+EE�}��ꏳ�W����"ֶ��2�BQ)��I� �	53d�"=:�P�:�� �ӡЄ��R�d �yw��
R�RǸ�Hu�LbΜ0�Vإ�I�;H=A�PUJiBD�QQ,7\$ܤX� -Qx��>���8G����YZ�F���̢R��	{WG?���e�2l@6E|�Ǉri�S�~�v�����*���R�;�ˊ��g��v�J(����_x��h3��� 75Js9n�h}x��Vn�C�n!�|���J�Ӳ�5�:f\������G �A38A�r|�ݝ�#��a���$x"Q^�|�~�:���I�h�M��UbgӼKrXF��+�Ƿ�=+�T��m����&�R�늤���F(�2�J� ى*j��"�
 ����,�p~/$�)��׌�ʭ [F�&��']��8�0���+a����O:i�����s�k��$��S����l"Ȋ �~�3�a�m� j�v�hm��)���)�^�� '<t}Ԍ��F�"ҳ�5o>�Q*����`���H���X��2� ��C�۽#�g�M�rM�HC%�Ef��Y�Q#E�r��w�E��XD�7�
�\Ҿ��p�N��b:%dz��T��z:Bȧ���5���mH�����<�'L.v�${�*�R2N��"s��Jj	��v�l�t�����(\���DN�5�d�1EԿ(��� �����اf@J�w���1f���e=�d��);�lr�\�Y4�Aw�мg�W|Q�<�������M�,)�Z�pq~�;D��;�"޲eذz�H�M�R���� �5��"b�Ը�� ���е/��Wz��H,KH�e��7GQ���I>>]�03�o����Bi񅋒a��Y5�f��VQj�����P��x�f�(�����B�˙K̆��Qe~�M�봥%��e�� ����mg��r�����ɮ��hq�RAGʺ��k
�1v�y�ukuv��ec��8H�2���.���1�ԶV�$�fm�L�f�OuP�.u�¥?`������ı�i���(v�~��������)TS�ǁ�\O/-f;�v������l�P�1$�,	U�DB �ժ�9m�ix�]���46>�1x���I��iph`S��cb��=4��0ˮ���ʴ�bW�=���݃M.f�&^Q��
�3�y�(�>�M��T����ЄH�e=�Q�̗*�8{w���vs�a�q �� ��o�LF���_��;V���R
�淟�;�h6�}�h��2�����U�sk���� 2@��N�(���
�jˌ��;z?����d��	4YB�p<����)�ј�j�q��iǙ����IS��Ot�v�g*'Y�hq A��u��[�)]���h��t�(��F�o�Q�i��FBh�AlN��z���ڀ�A��ų�~�rA�!8vr�^*(UE���b���}_�z$;#��<%��qH�tf&�U{C����Q��g�� ��ē���?���[�5���-ypR#�}� �g"��5��F�`�����w�cy�N��7�G	v��&y4��c�x�8
1��g��� �-��"
���#�-�y�0�v�fD5����J�/,��XO�ӥف�/��c�i�3��)�b�]��wjۏcB�^�fG����֧�]D�Բ��6��n���;�Dyڭ��O)�;X�ux�}��1�Vtx�ż�Lg�}P�19t���)�D�u/� J�x�*%��D�$��`7�g�6a�g�.�f�rh�DϏ%J��=n%rکHH
�\�^%����O���a��>ֶ͓��c�r1{��TQ�ѻH��lc��P��5�R<,CB��+J��N��ꗿ�6%�v���]��׎�o�٥�����s���HY��ω�J�T��)L��ڲC͐�|��t�qgu�tu�X�V���GF(Zo�@K`��2�Еk� �K̹1��]�0E���"u�'��C���C���͕��'o�f�ڴ5B����tV=�Kl�R'���0d��(n���+#d;��߻U������`��ͬ��e4�V��O~`��vU]G������RI���C;4wQ�4b{�s�������6�A^��"�!�i�Y��A����nO��&�[��	W@����e	�Lկ�I�-����s�V;Ƈ+�}#���&J/�]Y���?���0P0�z���`,�����z{ld��ZUd�llE��ݨ,8�ۮ#`�19/X:C#_1�s/���]�0�üs��&9��$������|=��cp���S�KD�,���{�G��H�^�Ge�<5���^K��!��3b��j��bg��)W�M���\�(�rOsy��ᵮ��2�t�2g��<Gpt9�>�Z�(C��k��zGxS�-
#�ǥm\��u����5�|���D�� ��o	D��0i�5��Ԝ'��+���'�Z�g\�)	 +3�H�qe+G�-�^5}rL0JX�%H���m;��MX�ġZ.B���"��^!����7fY�� i�3d�tt#����q$AT�ϥ�$ؾ8�ɆC�}�]��ު^~�����pZ"Jx`���l��aa��ST�ɫ�i�SQ�۠t���(l'�~!�(j����wr�́\͡vM����m^Mߨ�Y�g���C7au�ulq-B�:�Nжh�S��i,���Xh�; v�\a�+hqZ�W�������� n-w[���PhV ]=�ւ�3@�í����Z�$��x̹��e��?n�Ӽe?��\EMx��q��!�ͨ��^� lΡנ�GVˀ1#eͳ��A����?9d�:��FF`)V�֮�H���<��-Y�^��W�-�ޢ��:T�ρX}��e?1^lJϙ����������
�5��C�[L�7 P�KcQV��DS�ܷ��<ִ�s<#�-�WM\���.nTR�}��r�:L-§�O���������?��^}��]D����ЖR@\ L}zD9��koR1�ϼa%�-�Q�����ј�L�ߚl=n��ő��p�Gɞ��Oj�bF��T��%�%\�\�mv�s.�.���L�V��a-΢1�~O���dS���B��L�̵�K#�1��䪅����'� ���@`��Lr��=ap]����'�g�П\�b�,�����A/M�*H�JĶ�y��{!섰�uu#m�^U¸n����6-�Y�+ھt�D%���i�r��kY��36���@ਪ!��\Z�k;݀چ&������5�A6q�\��pW֍օ±>�_Ƣ��u����.��Դ��:�'� ����	���"��1��9��	�g���"DsR�1.�Nj��p�f�P �@�Y��E�y{T�?�Ad��f����`\_�}�Ob�F��h�>���;�u�8��I^��!@��~���{��a��H4H�5g�xe���3&�-���R�f�ə���5������Ku�'�������!],Ϸ�ʩ|�a�`50�Y�~�0�{�Ot���y��τ#��
)�� R܆�7ւ���~�%��9)��m�@����n7Bxφ!4N�,�]�8d��M�K>c�D�w�\l�X��(�w�q$���񈳮���X��E���(+-���A0�s��q`��<*K6RF�=wx������g'��b��y�6u�Z��ћ�֩T����ni8+��+�x�)CI��b�	j�Jq�M`�~>-K��9�KX ��N;;i#�x#�i�4FQZ��VA91 �?��,C)o�#�V����} fU����xm�hk��m��y�7�H�7XA�m�bp'q�V�+]sKslJ���Y6g�e�C�\�%���5�.��0]�����]�g�"3Y�l|����6���9ya��g�P:��bM��i�����oCZÑ��@ǫz߹�d��=���(�����_t��*D����`+3�9��^>$�����tN����i������dzq?0������r��Й�H+U<�%�y��8���"�}�����n���H(�ː��5�st�,��+�dD�;��������V�5���'ݱ���hm�q��8�&-��^����]�(�f��E�;���]d&�xٟ��?���p.�v����W�9/���i���c:�.�^��x#G�	���NԹ8[��E�k�[���,f��ʋ��a��|%^G#�F9k(7��}nosVD��!۲"��N#��q�){ss��	S �1@D�J�+�j���,��Ƿ��qN~�Ӗ�$K6S���{vk����pC˧OX]M�ǯ��ȽVب�!�^lZo�2��Ξjȅ�>�e�������{?����l���S��"�`�>�H}4qɩ�a��&x�°�Gk���c��˹}����fu[Ѧ�!��0�i��>d��'B���Kc�g�s��߫� FK�tb���;H;[���l���
o���h���YO�����{~��� Pp�9��3�dE�5B�S�ڹ�p�[�]�B#t��+m ���^�}h�h��;B�+�����=~M6��<�����~p�Q�_�e;T�${�@���!�'�#����e��eB��"�KG+~mĀ�#�������	�Z��ݯ�(Ö�b�'��Q:��L����b��^�b41E��1��� �T��a���c�t�l�?�?���^6�^�!L�D��xM;���b�	:6)�vf X^C�G�oK	�-)��V���s�%-���:���"�X�5�:遛B�`#j���v<��BR��f��Xa�Cȵh�:��e疣BV@��-��}�q5d�C%����u�?�,?�2�a�O�iͻ_�2��[wLb�,�0�J�R��B~Ћ���:[�]���JX�s?�zx�*��S2�Y,qu�Lc�!��q^��������o2�p��Pդujq�@�I���@��@u(�^�=�6{q����O����dbj�l�<#�/©ڃ~$>Q"����Ć0K`�qƓ>�I�h�U_Q��K��u�O�"˙����i��
͏'�8)�<?J���累�k�ow�!��kߊ�?�JU|KD��!�(�����.2]�3ڈ���>Lr~u z!��^�M~�D��uw�by��R����i'xY�[�l��O��a>ׇ�8=�eY(��f�]F��ᇥ� ��!em:K��|#AC��*��0q��X������	l4xH�����oCL�mg)�}���AjO����"VN>�Gn��(�e�5�pHZT�t��띷�EW۶�w�0�ǚ'������f$F!�<��MU��͂�$�;r���U�H�,���̼Ti*��M�,<S�� ����ד���m�gcɨ���/ִ)#�Â{�Ƕ�b�C���2�W��!\��7ǉ��c�d�_��\�T|�e�zh��G�}�E��t�:�$Gt��j�9�����
)]pM�E;�*N�p�v0�
�U�$�@��FuԗN�b$ӡ}�PN0딟�O��h	B�2g�s$W U�R0:����5��h{B���ӗ"���Q�do�
���u�G� ��+!�r����8���'�g.H�g�-�`V0�.�6>��W�7��UҼ��搅��`V�qq(#l#�y|M��K ��<f�Z֢CtA98�f'�6ъ�vC�1���baz��j�-��˺@4�ݛ����4D�=ǩ-\�
E����Nz��K�O|�9�?�5l	�{��EM��SG��!c��nx��{E�h�a�\]���~���@��@l�Ͼe��^nM�`i�{�����VO y���O�󬈒���1��r���%�a'�v���b��}���D|;3;�#��"�e򆑄���ֈY�G�����Ǹ��)	�A� �*PiY�M�mc�1����~�����A+p���}���6��u�@t-3�����H� �J�)o�\��ǯBS��A�b��
D��ͽ�+���If�_����_K�ȷ+i��R����S�M�V&����5R1=�߾���,�uH5��o�jt.��M��o+���)KP�)2$�6����ar]`\ki��vCr�W���]C�Yu�J!$�|T:|�s^�蟃�GZ��:�I8��+��Y�KŰ2�&j*ԁ|�'�8�pv�E���F��Ɂ�؍#�H���.uqr�-6�L���~�@�Pr�D�{��xC�}�֏c܃8K�i���"`s*�~��
��� ���B�A9��w��ꜧh�5���NJ���XM�T�B>;��눮Y�8P��RZ���I��&���\r��mQ�+��Ȥƍ�y�S��� �p�⮠ ��!�ֆ�8�|E�y�D�rj�D������A�v�$�|�Z5��G��*��8�pu.�Y]�����n�*J~��Һz>~�R�K;r�8c)�0MY����a��SF0�>�B7u�6M� j;��*ɺ�F|(�L^ڥ�=��'��_�wnB@��UŹ�b���Ar}��e���y��/�ĩ#��z^�ϖ4�M�B�뵼%@DF�x*��}��Ю���~�3hL��E�>L�������M�c�|�9N� �k0������/���Tu&T/Fp��	��n=3v�A�Wq:�18��7PH�[}ɻ��t���'rr��Fc�2�	gz��r0ѣ:Y��,���e�����w��� s:@�&��R�h��1����[��hŖ���j1�`����"4O�J�
-t8�L�ӄ�����Kk[��M�r��}*�mH�1Q��DWBF��~�(�C��t��E��Bj� |���ʥ	PJ^�.r;gxvw_B�߸,�9�����N�c4:�O]'�N8�kx�2�9�t�kc���r���בOj�ɋ&l���V^V4�a�H�xF�kG7�Et��H���jm1ً"�l���f{j˔r���B1��-u����`�z$��YL� ��g�'/ga*�L�����Σ�۫7���B QT>��A��01Y[���PVew���,�I<XR���vv��.ďGC(>J!�[ƕ�V�y}���Ŧ+9�oM��ۿ! N{��,y��&�EVB���������A"�N�v�_�{m��BH�O��!��9U���.����n�w�TB��A��2�U<�-�� Ny9W0"*(Q�x�[�"!�x0���W8C��eut׺��f?9T���*���+
k��lWc�9G�߼���]Hy2a�%Ģ¿8��0��	{X�a5��RQۉ�j�хQP~�/R���_����B��e0@�Dp���+ �*1˶
UF�ŗ���������a~�&^da"�N^Dq�;jq@�pkڌ�'���uÂWU	u��=���~�5��N5}�p�1q������b#���"���@��	򾏡]�����'YOOczWJdJS9Q<s���i�[�ҩd_kݖN��rՎ��O�v����q+vd����������	
~�Z&kR��;�"cbn���+� b�v�Q�Ŏ�/^d�B���6mf��' ���p|z��|wo�Z���pIo�sܱ��g��+�95�s�8_d|�����6�� ����{_ZX��6Yj�p"��!���]���{$Zel�|�,��!р����X�qך?����ĞOa(�G:�7��)�>��v�x���S5Q��*,?��Q��c��I"��ѥ��c%�)�V�HM�;�X�:��t�O�O1Yt:�Ӄ�szG���g�L��+�'k6�56�
�Y0��C%�d��?���"Q}���a���@��@�f��?�~e�W�ʠ�|R�⚷���}��������`���}6`��p�[�j_���Yr�h-� c�D�5[o�m��`�R��xc-2mad2�q*��ۦ	��ꔒ�R2E!��;Yp��_5L��+
d�dR0��}���1L#;�~o8|(��ƴܲ�
|W��B��Z��O&[r�5��
k�����%DE#&>���}�����c91(�K�71p �����4�G�|&�L��F8j?l7���y{g|Ӈ�]��<��<G�-���6f�O���}a�|@����2�?��C	%�j�V�ui�VG� �s�	�P=J"�+�*֕�Oh�ȍ_o"��mݬ��eOf��M����)��D�B>r��;�?f����(sD���Fg-1Q��p�0�-rԿ�D쭭��4m� ��a�K��Ɠ�me#C�m��[�	ζ���yihp`&�S%�J���X�a\���ޏn�#Y +��h���g���Ѥ�*��T󥥑�A�bO���	�\��P_J��	k:���@��lX5w�#9��4F��~�e��y��ޘ+ĸ�1�&">�����g'&2�$���n���Y��庬^����7̾���|(9Mѝ��?��y c�\Kj��*y�-[�v��+j��,���[��S{�g�����>����P������%�'�0�n)��Q߂������� )�$�$���I1��;����X4A��Gt_/���W�/��<lt��ክ��?0/N��9a�_L�*�p��I&��&	�3�}��?T��#v�b�y��[��7<uM6[⯬x*����ƵD�$����7���s�Is�a��8��u���#�!�G�4�%���0_�bwpc�I}�T�aL�E~�ٵ�sB4|�ηJ�#?��v�-�[�2��<5�U�cH�݇�� S���r}�ܦ	�W���4���f:���'�)�hZ���f�k���cC�w$���4�iAu�#�}QU&�t��Z2?����i���b%��M3���C�d8i4m��]��g�
�P�!+�Wf�̙����R���
i �/N��,(�CIYW\�,O�_�g�tp>���2v�[��!e2&�0���rJ��kC.���s{�����+L'F__a�O��7�W����q�.��Vh����y��
�����F�`%�c����"ac�۱�şO(��+�<�|:��3�s��%�N�+�j�YtTy��f�|8қ�A��ሕ�*�n���:�rF���'���)�8���n
�M���!F���XDD`�n�̘��f�I�A2�q1_�o���:*y������b�~�;�� �~��x%�)�t��rg���	�a ��Sl#Yp��=mF��4:�]��g��NFs�_��0zH��	�C�:�A���)�Y��r�H�^���NZ���Y�}���1�3N�Y��X>�hu'����!�Qd��>j�&J��I�}Zf�k!k_�UU�	��4�I�r+�2�� �$�Q��j��i�Vl�tϡV��"k}��ژ='#�����/�^�f
vY���':~G��%��]���>Np���szj��%Y�8��t@�dm���ѷJ�r���c`�n��P�Ψ�\C^����T,2��!� �]7oP0_&h��w�>�9��󘜮u_E��@'c�����K����\�sX�K��@v{1r�iV�l�Vo m�
������0FK��@ `�p�u����%[x�!)�*&i<רMø7_��a�t��[xX��R�:��Nzm ��.?���7��h�Fr�,�B3s���d�C�6���$I��JJ�4��wp��=�����1���N��>���iu�H��,r���Xz:�ͨ7m��Is8�x��桃]ږ���
�����H]ԭ��5+��b���b�mP��JO�A2�����1C�3*��=˺�ՁF�0��C��{,"�����Yi�"��F�ްEu�h>�=E��ܡ9(<��$�C(���R2;*��H�9���[q��N-�(�=b
{_�o܇ا���sh��~y�D7���0��E����c�3߰��eZi�$[�_�����Ju�v�{���t#�u�) ���ސ�	,���Xj�0�v缪,�b1�2�s6'!�g �S��7�E+|���+�fT(�G^}I��T��2��W�r6�MB"Y��Fz�J׊t���J���Ǘ�mL���4��7���x�߲)���jK�p ���UF����	�z"����[�谒������+pr�� >&ʦ�abp���8��L ���f��cMr�#r��D��G ����zt1ej��!c�]|`.����#�a׀8��KDL}s39�Ʈ�A�S����|���2$]��s-�\�y�D����W ���!��9�@�H8�O��LU��'�!>9\��31��t|�Z��2_/�@�l��Nr�k�@B[1��u[�	y�D�8Ny_�Bfc�j1�ű��x�sMA���}_Y���H+�Y�\t���k���gV�	����y���bٗxo8ap
M�˝�Kbm��
�0�!o��K��2j��h�/W��ӫp��|6G�m��Et���y΀9�̶U`����Q}@�-{�!��^���B�N(��˥D�� y/�fd��'xw�X+��Z�O01����z�������H�KY�� /d���:����C�w�]Sx��+����3��I�Fh�dΠ�%:����o �.g���7?)�#�g�=Lx�[��KX�/b���c�ۥ��'����:���4�x�>x�1�@��&0Cs�u��ԏ`H3��n3�*̫[��a}Ղ��WǞ;����DLFl�G~Y}��	��*�����\��;�������9|�����&x�`��}�XY�C����1�h	'���ت������(�k��u�`Z�Y	�1�9�Ly�c�T��Yz�(Va}�ɲ�j(�IB�>|�>�����x�>ATA�r��3˰�H��.�9�3��� ��I��c2��Z� X| :�01n� ~d��KZ��á�lZ �3:t)4�Vd�[L�B���j��\������sj��"��1��V�1���	�_�P�7D��W�)��th'-�أ�L����%HJ��r�uM���.��D;�~C�a�{��A��*���+j�{^�YR�i���e�W�z���c�P;������/Tl�l>Q�F�b�0ΊJ����%��}��z�Q��Q�3���s*��g��d*]].8L���zS�cҞ|�_�/��k}��H�P�Ϣ�O����/ ~�2�i��`u[*j��rb/��g�z��f�e�*���E�;��U��l���g8<�U%n���@׋��4$��y������4����Ҭ۵�"�;؎���|��.��'�L����@�ߘ��٫H �/"nu%���@W��bX��B$��K�|?��[�0���&O���؆�D%Xị�ձǐ���{'*V����
��!,�2��j�k#�f�j�6:A�歙���zf9q�=��K��9��i
��z�y���fğ��5���+(���!HO��q�A�������uQ>��L�H��_H�
üj������t��Yn%8m1��3j�Y�c�{�!�鏷bY��j5���J�k�Z�_yz���\&+|��<�Y��̠(Â�!�uI��`3���$��= ��˂�8�+��X�t�btD��%M�+�(D�fI��im3�I����v��(Ly
�C�H~�\ݍ�W��B��%�nu��B�t�m�+x
QN:{ͯJ�r 5�w���VH��2a��� ��u�Q�̇̷cN�&,�U�(R'�n�⡴[J4ZZ��y���~�2���乪|v�F��f/����*e�=��|�'�w�QP�F�����7�+��R��\˨Ґ��5��V��1�8���1sy�e·�x��Xy����hR�<Sη�����uAߨ�2�t8����tx���EJ�۞	!o��])l�6W� ��g �_����56�o�C^ө��^
����ER�,�Y_�/<�U�zj���E��<6쵓L��&�s�K���L��a�Ƥ,�����QP�3�P ��U�6�\Д�~�KO��5J"�q��VxE��'��ɞ�NG�Qm������`~����2Z㘧��88ߜ��F1�R��"�LNE��.��U�ع�nv-vM\>*)~8��t�(�l���}���Lv���/�d��E�}��S���P�/����+�R{d߬2�K7O��eB�
(5���YEBEj��(�/��4��(6�T�2A8�6ߡ A�a]��N8d*�����%�Fz��t$�7�u��;������EW�ua@�ϳ҂�y�>���L�ma�q$�U`��z��X))ʉs��Nʗ�L����"_`moS
���4*~V�A7�]�x������ts��N�BA��
-n��,��1	L�Tn���Kו�Ε+�3��� s���-Xr�(0B����������єDD�C㹞G��@�g��!��[�p��o�2I�32�I���,>��y�0Hԓ��i��}k~�}��������b�?9�v1<&U蚭=�1�����s�.�x2N��x��%��4b@�(E�&W^ﭻ�b��]��J�W�.X�#P_����5�mN5r�?��s��b��!a?��rO ��PV`���Դ�
'_\5D�2��.���QG�q��ʱ@o��N�'H�"͚E]�7mSqe�;�gw�,�Q��@�[�UF�W\�)�`�ޥ���M�3�����;b{]%S�#��v������j�٫�Q���a��r�t�{K��7~�����v	WN,��|0�*�$��½���$����f��˸&޳�y���*G;=���$�Hb��c�}J��N��`���`�\]�̶�K�6 P���*�Vh<�w��Q�Z`&oD�8R'��� %~4�P<��o�%t��[솲��Gm9�!����L��@���H`��V��KcE��8B�#�on�હ�-�˹N�m�v ��:˲EÛ%<���`a"���������~��PYr˺��|)���x�$��I�p��4�K�ˌ A?X�K�4������R������?#�|�&������[Yg�F�#[�3���΋D��B�����7�j�� �s����C��֒,l?n�����t9�]��� χ�2Ej��|�h��@�����k�Ll��n�OΦ-�����}(���}�Z�N6�II��e��e&�Ĭ �{�}?n�Lʀ\����j ��
*+GowM?k+O&�1!!π8�!h�$h�ۈ@EsU��	�%�f����1��d�%�+_PU�kܖ0d�:���p�	�k�<���/9��0�iA��:x����T�+=ˌ�
F0�gILh�N;��^1�b�8�N�s~e���Ѷ�:�Z��`�i8��� 4�A�=�]oy����K�a��#l�9&� $���ݨx�4����dJc{�~Z�_�S�	?��F��ىB��%�p�{�q�R�)��㬺n��/ xv!�R5�Fƻ�β�g�YU��81�X(���gY� ���ک��>h:�,�`s7,�����b8��Py�t|�Y�7�3.H��k�I���f<�{p�g`�ZM��5�8ޭ&��hlwbNY�-�C�[L#��}uJ�ڢ���������N򧌔�x^�M��Lͯ�9!�T���W'�5xą��#�^�>\��@wㅖ����U���*hޘ8��Z�U ���$�Z�"�l��u��9͠6���F��}�j(���6;6}e֔hc^��G�I���j�M�Tq��O��|h~A0�\H!�0�����mP���I�g�ލ�Hxw�+�Ԯ�
q<�bln%?�������(o�%Ag$Csb��B�ZT�I +����6!���5ZPL�q���X2��5+`��nn#���'X��dt]�?Z��'�G���yPD�owr�U^"��L!JO�#?|u��%)B&�c�_À}q�[|�nK�b7�F���oJ��*���P-.��;�+�BG���=��+d8sSq�&�.���6��`��a��iӁ
/#��Iߙk�:�[�ђ�5��R�I	kqMVc&J��'���Y~�R9�<��T]0�ľs�n�ۊ�ƺ�T>:y)ձ�4��Fa���q�?��q�/��|F��.�r� �rc����܁~�]Etp��vOK�����n��+������S[�%.%ΌU\��`�jz
:O{q�^;|#�lh����0�<�=��g+�
���VwD�8bH%��zZ��ّI�'~�9V��<T��t!b���U�^�>ef����U�U~a��sJ*���(�^dj���CG�>ghB�Ku�]�GnP��]E0$#:oz�(��\˦_�ʅ�����O��SV�i�_��i��0�2�B�R�����]j�s��bl��wU�(�q��֧S(���H>*!������P��:S��W2��������1D�ŴO�^>+��Tj�%n �.�t����=��w~���� XLNo���2|�y)��S�y�r��i`��ׁ�\2��@ּ��[�����n�z���ȣ�c��^m}�b�����.�w���z����<�$��Yװ���\=]��a��X���bS�)���^����/h���ʀC,�mQ��#�6��0����p���g-�6�D�u?U�9�hP��N���J�	�;}6B"���bQՙ
�`8ʽIP��V]��  ��U�2�,��F�TRfE��������)��0j`�RZ��>=oq-���)��aW�t���s2��̑�������10>�������9E�ߙ�c��P�]5��!�k��wx+AF�.Y�X$h���x�皣��W�$9�Q�&U :`}�yFI��&g�
͉��s� ��I�i_]��[��uG�Н6/�o.�`�nNz���k'�D�x? 3�2�|�lG�zT��a�«w�?̀Y����{\�-�a꬚B#���J��= ԛO�NEu�k�I�x���s��Q�������
FEB��V��^�����	���~��"c�"ؖ��Az*�7�W*����Z%��ɶ³W�6RQfp�i�F��q����|�7�I����N C�6�9g����#6������ڪ`�3G!l�x/ޱ��?�0J��͂�M5*�����U���%`(���[�h�!B���#�6;�ps�o��h`�r�D~��S(�W^�'و˨Lvm:�7f���_7�}p���q����9�ӜpZ��T�s���b���-����U`�8�'vW�gm�+}����D+O���#�1�.Q��A1��o%����M���Sp��M��|�ъ�2CS`d'u2�O���.�����z`�������_Z9�7l�M��[��
��:��{*S��f "( %h ������Y�w��Y����jM+�i�e���A������	>����5)Vt���j20��yT��4�ؚ�E�a�L���fZl������u/�*�w��R#L\�-ͳĕ�y�F��F#��'/q1V�J��J@꿃\R�Ϸ����h����7��ލ���U�O����^����rr�tRE*�!�� 	�/N���=�c}�:�Uɯd g���߶�o�c��b����F8\+���	�-���Ac4HD0)\V�>opye���4�K+��44��u�Ş��^S�<��;E�=ʇ�K�%��ѹWرD�������HT�j��PF�ӭBjeL��j��<'�m�d���9)V���m�z�蕏D3�eBC�q�H����-�%�w�
�`,�u��H��>�(]u���]���䴵eo�DBH�V�H4r{>���2Yx��F��'r��%`����]?�R%<{��2��Y�S��}��Y��Y~�Fl�،�
1��U���_�*�}�~@9$��)4��M[���K�\6P`r.�W�jd\1�b+MJ���Ŗ����Ɏg�#�do��#�&�Z.B�؍QH�n��Ÿ����c�,�vm�����5;�1��X�g�u���`�S�5�dز�KG�j�"7��7Y 8_ڴ�Ȩn������Z�S�T$�c˰R�m\�DֿL�	i��4�:ku���]IHp���?�n"I��}��բ���(b�ųnǝVZ�a�+/�,�8ui�r��b��2r�������&���g@��p��F�%��.�������[;�3������>fCR&P���I�*s���VxW�%��d����w7���t�v�7NUN�p��4�<�?��$�p�2#��^�z!����s/̀����uy�
k�o��.�w��dߕ�����thP��'Z�0�20����W�o����6�o��|^��g�ͬ���b�N�,��Bs6�۷(6�w'��h��_|�F�����W
å~��<����툆����Z����mvߌ����w?@&L��ECT���Ɖ�F�Pp�:c��ߗ�L���;;��6 �쟿إ�A�Uv���5ŀ��ʐ��|�SM����FR{79��Z]G6g�����s�E�	�U�q\�������lB��,7��(GC1�<�������.W����wpG�e�[�Z�:LZG��ѯW����o���6'D4?默�D�d�P��)�Oi߱���r\���5(�E�C�Ip>�_|͡��O��o#cˬ}��$�xB�r�����^���EJ  Z��u7�3
�
!4ay)Ba�h��v�۞X�����4�:���0�����Y���[��,�̀�����r?�|,3�'y[��):wz�	��Z����ǋ�3ʩ��W^���\wW9���_o2��&�h��ʊڬ�7���ڱ�Qb.6gL&�q�cd/��	��F�f&.g�8�-����9L=�$��T��E;��[�zydM��/�K&<v�A�x��O�����D0���/ͪԤ]Y�},�y�ff�-Fa4䵞���È��~8�;qO��>b[K���i�5���8��%=vIl0��Ϊ�T�(�oѾ�+��iO�"�a����+Y6��2��Ϭ��?Q%z$�i�/�c�)��g����;��<��3Ӏ�ҦAj�� #qaOU.I��kJn\�m��,�Kf䪻 ���^,a݂�:s{ׇ�6��
��U�녲KL�|C��-3���դek�]��lQ��r8�!&�ڮ�$��������du�'D�p
��o�.��G��o��6����x��:�(�Z�'�Ek�>g|u���� dN��<"ܐ/��Z󉞎4ەGvڞ�b��8�0F����	�5�f�E[攽N���/��AS�Ը�d����ʶ�4�4��r³��I:Je�\��E�A�q�R��=���f.��c��C� �(��' �\��ꚸ�LeP���T��p�<�f�kyY���+2�ۧ�Y��|����`/��k�Cl�d�Br9�J�Csq���BXc�Q�F8io�4�@����c��t|--�K3��{K��e�~C�W=���r��/W-Xz�J����Vƶ���}�=vrgg�J�x�K�Y���oTE�f����Pa�QA�L�xM	'jQN�%�g�+J�(K��g��gG����>�~饣M!�F�xaHg�}�2I���V�����J�-��O�qF�#��2Й9��~����o��u�p��~�o�MȘ��SJ�`����)5�ED�o7f�gE�=���"��2�����;���ɑ�6[��k�z�˯Ƶ�H�������$ŋγ��@K�Զ���Q�[8@<��/�VjKĔ�mFa���W"��P��O`}؊|��Շ��b$n���N��1;�Vv|��;Q��+������$�Cͷ,��6X��_���B�_�/�M��>�i�A�R�?2Fu9��c�A�Y
�[:H@i%�x�Z�������c�g����f	�逤j�y�M��y'�	'�9����qtr+b��?��t��/�ZSw��N=2�fR�I��M�I�"�ap< r]3��������$k	0n��-w0����}v�k
�0^LM�n0'��;P�J��a-���HAT��S��@�i��M��έ-�G|��ҋ�G�
��k�2~�1�O���0 4w������^�=��V�r<&\{�ϫ����:����⎓��!R{�_�Sp!j+�&�\>x�l{8! ��)��ѽ���\��&��p"KoL��'�B��	�e�K���_��oU��H�T��SZ��\w�S�}���i��7a��~��#������ʤ���tY��W�[��]� ާ~�-Ynȕ��N�Լ�W8������q���^�B��w��:�d�C��qSd$��i��+>����3TV7�D����K2�z����aⶔ~?/|�C�����l��su��S��4����D��f�Y8�n?DNlaN��j�ǖ����] Փ��>��+8m~epR��`�������pB�0�\�A���ɡ1п(����olm,���RKBJe�TJ�8w	[��2K���2/[�eX#��HF]�>6�
����e-�kEf�!fSZ���GB�<�9����ǜ:�D1�K��C��N ��e�G��Xa�~�I���"F�D�},#]��J�t������㬖2�����$|v������ˁ\|��VVz16[b)�y�Bj^n�Xտ��+�6v��B�X�<�
|��S��\054 E��'k-!ȃ��u c>X�s�y�H���D�Ө����?5?{~Z�r\b��li�*4~P��t[y/,��]�"�!_����¹0��0����T��).�a��6(�х�Z��	�����2���`��@f����O�ף�IgʓmҜ^��:�6���dNk7퉈��ͯm�=$l�&)�w���F!�sI�)gs�sì�V Q��Zc��))�ov��M@�����vxL�ף8&��d����3Z����Ke�=}���]�܂��|z�]����ku0�4ݓ�9K�����>�#��C�S�x���u��a�6H<�]r��M@��i�VѣP��@�Y���.�_��Y���21�]g�\ 2mM�D��_��0�K�pKS�����}`�7ne�g����~K�$��s��[��+�׸X��z�jWؿ%�3O�Ú����J��y�n���Ǉ>I�߶�3�n���VV�^5!q������Q>Z��� (��,D����3"Ӣe�^8�o���<�\)�p��0�(ে.��m6�^�X���)��.~���2)�<��_�k_����y'�c:�q}�<#(�B��IP�+^��
V�w�T"�va��pM�f)U9V]f�!��S��St�c����Wp,.l�ȳ�Sg{;�+���$Hh�>Å��=a�Y�5��9U�β?�����Q����b5
��y{^�*��؟�<�9+��1�sR'���i�g���'�
6��x4�՛�5�r
�z.�
�) ._@���\��{�3��IY���rD�T3�*x��^ �f�ϕ7�5�ʚ�<n̙���D@��!��c�\ѱ�!ޖ#�y�0���P_����";�ʽ���Y�@�M�R�7�J̗��{-����l�;V�
��"��F_P��.ToaM�/����3�B��a]��6v�|�/N񨵖�`C=YA��Ā�{�����,_Q�IYw�����I�hgLH��e���

@��f���0I��$QC��xD�F��)��/Ǫ���&ʚ���J+�τ�L\� l7��*��;�!����@�{��J� N�fòTbX�]ܞ�W����HXq�a{��qL`�_c�cYJ˨�J���Y�"`P��C���]��C��Ӡ^��)�ۡX���&_�f�D�ǽ���<�o3ū3�Bw`I��59x3�$;0%j~!>�A.T00T�tx�����\��D���<�����ti��{~m��襝U��\������87���8��7�ʀK���s�����<��1��3�W�ו���s�VK5��Eޔ�=ro.���X��)���95d���v�r�ʐ�華�$�3�M�)����irQ�%���g�m�y�Ł�?���}l�R�F�F=��k�� 6��X�Q�P�l��Z��S��Wefg�[��]���5[(͒;q�^`�ndq�K��:�Gla��!k�N�iG�8'��P���YD���^�>:9�4��W}g��5����&�6Ax�5`~0^�xzuў,ۦ�Z�#�
�!B��,�rݙ���s��*�B��~��*���!�w�����^u_�{�5�XY����[C̢�0�<<���F��B��������Υ�[��0��{��������W�Bh@U�_��P�g*瓂Rc@�A]�*�A�%|1x�<��,i0?����8�3��i��U�h��K��FD�p��ꋧ�����K��F}G��Nj����Dsy���q�by����Obqy��f�%��/�)���u�ꩨY�H7�x꿳�)�����H�z`J�,��錜��˧h��,�n��T�j�M�iN)"l�?ƭ�c��V�Ce�Jba�oGk7
�_+hE�2����!��v�3q�䳳����(4�4��5oȅ ��=���W�|��ة�˻&��r�+������P�ћ	���xe��a)R!,�6���#< ��)���E_�y<�8[�˳�E��m�^Ŀ�Y(tެѬ	_H�DP���ML)���v5��YV�	����V�6�W��o=��	�Y���]�{��$�H	�ʏ�3 u���B	���xn'�ui����k�!�1��J'V�_�/ݦ�h�v�����*���4H@�=b��y�4"�@�گ�U*�> �7��Fή6h��ґ �-!��f���h�zb��,�����k!qOS5i�_�qW���}�v+�]|GG.B=hViY���z����>&$�	1^��OY�[P�;?`�a�09�6/q-�n$�]��-���jD)�*�g���Z�b�PT�s%�Ǹ��
�ڂ��[���F��ջ��y��o���9��(O�҅)�� �����8Aȫ�;g'���s�����*a�
�	�Ts<|��c��uN�mh?���ku-˒X_60�9���R��I{�f��F��L�~�h�]�+��.c��rBZ;?r�f�����]��P>b];�f��U���|����ź��i;��ly0zS9��ч��v��	ϳĴUO!�r�cP���	���=?�N�X'Q�n?Q)@��@|r�� {DJ죿�7��p6��,g�*�i���Wʓ��1v:���/j�"�z��z��:�ke��h{،S�H��5Mjd����ts�sc;��i%=�D��ޗ�$����Q,�:~�ªM�p>���	̲�k��ˎ6�T>ѕǆ���4@t ���w7TC�j�1��k�
����=�2
�S�<�,���_	�`l��g���R�0"�8,hӳ��6e�%�R���ؑ�1��z��%��'��?T��5�X�|v�T��D�}���+�7`ě����E�N��PǸ!�U�és�۴i�II���x�,s��=�*3� ������{`@m�g<�� Z��*��e%g�4x#s�{���6�Vj^��M���#X��m@��o���,]���[*̸��6[w�\�4B�	�~�V��'�9�JR�YW�4s7Xm1+ޝ����~���ƦY��q�F�'�W݋Q!W)�
ݟe���>�ޫ
dI� �޶�HE(s���*�
C_�L����P{Đ+g�v�t�V�f'���Qk"	O�T�Cx�jG�ea����8%�"G�^?E$f���ٶ��ꅞcTb�lN��Vfq�X��3t�_J�x�Kʚ:��{�}>����n�t��̳Q�{EB�\j�%����/��Ō� �x�gz	 ��bG�1�N=�9�o�}� ��ZHS�`�\��T2@*k>��0ſ??k��^��N�9�u���L�X=�p�SC{�m�L������6%!�<Os���k�I�9�sq�������sѝ鱚���y�Y<��w~+�HϲEu1�T��� ���(�L�胂�Up��Yv����LH�d��$�p8�=9����ܧ��lx'���܋�o8F8	��U���lb�{����.r�i
�|���j��$.�O��T�Q�B		�1��zq�����Ŋ���ڄ� h4����p��D!l�!���,���ئ�:,[�Z����y��s&\���_7ٚ�d���n�=�@�Ҟ����M�"´�"Qc��,]�����^vZ�#�pV�\�33���szK�6���@n,��Ë&pt�-Q��W�cą!Z��F���Ò��9+����?�ܱ4� �D
!ja�e/؋�8��˪�k�V�+��)����
Wɪ�fJaQf�����H��%9[@\�����?[Sf���������]iV̳J�7w&�W������iA"��zz������V_*L�9��j��Q��A��$�0 ׶���$u����0(9��_D��g����}���	��YE�{�Q�-�
%W2�ȥ�r+ޙ�C��R���	CRc'����S������h�\R*���ܭ ~!AF�wS,��֋��5G�-2W9��3�rܡ���.ĕ�E�:���~���R�������
jb5XE���8�8󂐃�{�`���;�j��֑]�[nf��p9s�Ig�TEW�N�����C��5��P]%�)�"4>�\/�ո��C�ZI�NS�����>j�t���$�:kP����M����=�K/sT�⟞�v��B�@�˃�Q��Ƃ@]R>��U��,X�"�=\�	^�A�ޔ'%�z�����n9��F�����"$��y�U��gĿ\��J��N�ᘕ�Z���d�f���q�mi�!����|C�f������;0��"�mF�Z�_y{�eUR�	n�x�O�ƘM˔�Rj�.ѯX��pQ0���BQ�����)l���'�b����Ykqָ���ǔG��R�_��G;��pkE��� ��F����|���應�������ھ���ʰ�o��m��Ί5���ָE\�����y��d+�V�]�0���R	���b����)[9(ȡ5��b ����u�3��ą�/c��7e�����wŴ�X���ɦ@X(�h9���������R6����0@\C%9��S�7YS@;�z��Ť��?��a�v̌�J��:��~�k�`��F�di�,����ߚ�KQC��!�g�����jv��
1c�P%1�_R�4�]L��ﾗ=�w�'��%'G��|S31�vCߡO�B1��a�M&���/�>���������H	�&]��a��&����,q_B;�`�!��_��U���c��JO���wZ�5�X�	-R>P/9�I��ӻ���8Z�|�ӱa����= _u�	��D�冺0ԙ�F/J*���=�Ğ���[٥�랪�YFy�#�z�rbo�;d���=�xk�՟�
�EQ�6p�)�����AĄG��0C���b���3+�$G���4�I#ZP�xґ]�����B邴��te<f:�]u�`�B{Boi�Ԫ���C���N㷺?m��������a���O�r!144�+4ŅT/�'o2/dy�!q^�����kc\�)hY��Q"-&ɤ� m��Y5ep��00	��>G����魬k-1���堊-�15y(�`u3�a�A��^b�O�����¾j��N'xg{Rڱ��M�|��G��^�sM5���9�ֹ�7��m��2��~[�GѪ�/V�.)��ȸ���cf�p�-Ӷ�C�<h�F�w��`�>��a�a=&%6f�ΐ��TW�m*����9)˞OHuXC�Py]x!��\��j=�mf��r%��Rh) #�5��~�kހI�m�a&��C�,��c��"��Qt� }Ǻ�O�,a�� aD��uo*��_U���V��h��2�2�[�$��[����$oF��#���\��p��kL��8���.1�ᚃCu
wp������.�٬/�h���D|�D_<�a�����!J�b^Kn������
v�b����.K�����e2�w'm��������)ۿC�����V�?/���>74���di�J�vzn����)R*'4�W>�;��J�ޱjl��2��*K��&ZpfV�ϪX$, �Feꚞ���L��ʘ���r��� �m��J���<@������M�z#����8C�p�;Le+�Qք3�em<�x�Up��(b=B`3���.i�r�i�v�;��C�-���v|��'D�:ȳֆ���ί���B�����?��jJ�P����:R$����fgB�Z$���-_�1�L@ӫ�C=v�Z�����W6�}��Zy_ν���������jQ�L�R1�۾�n��.Ʊ�b9>�_y�|�f|����}y|��o
eerv l =ƀ�[2�J��j��y�	z�i������T������{��y23�u�xS����뱬hA��"0i%=�z]�>Һ��¼�89LR��o�c!�:͞��\�X��e䎎:��f�,���B�I+�oRE���	ެ%{~��"��ԣ�a$�_2�*q��#]����ؤ`��V�-z&�?����+Z���r�*9��_D=}���O�_o��Y�6JЬ�Q,��{_O@ �LW+�*3o��7Uj��#�:^x���}*���c3�r��Τ;��8�<����l����Tz����#f }�>_hfz!���%g��7dmS1�����KI4�>7�F�I9pX���OL�q�K���Gʩ � jl��2o���������w�b���,Ja���#�.`��m�B��x�/I�k/�"�,���	�~7�k�K��}~�R�{A�ة�?Q0�s�Wj�%��;��N��m�`{5�S�7�z�?T/k��ub�jAY0�z�û��b7���m�5�*Ƕ��'�*��jp'�٣
5rH-��\���1�֥.�����(HϹWX�=Ҙ�e�rT�E	�|TӷO�	�Cta����)NYY��a��ЀF wҨG�j�ū� ?0�P?n�v`���4�p##v�Ք��坁0D�܁@A� �$�]v ��Q��׎<��_���Y�/���)��:�%����P����3sx��c�n��Z�c��Y��]D�)9s����5���ƍ݁�}�F�����,3�q��'�ӝۃ<|�1�4-i�̥C��V�r�D�A>����B���gCo�k���U�X*�9k�D��jX��*Տ���Cl�A$��	aM)
�?;c3�`h���Y����ǝ� ��o]q�r���$\=`'(J*���5�������$�C��C���-�s��K��<�;9���;>��u����3	�A3��&��E8`�t�3�Z�ܰI�xչIf#���@m2����5��6_B�pv�,�E��Ǌ����I�
E��S#���] �TG�R��E�2���NM`����F3�'p�AF&�F*U閬Gt�|f���H-��)�G�]�	��nJ?@�D�dR�=ʚ�t5��$�ؑ�C�_ɀ�jI��SE�b�?��v�)�<�%��l��[C���f7f��a4;W�	y3�[++l护u=����A��I2>��F�V��l�N�Z�y�|n^��5�#�<�/���V��-nN�$�+��9���E�6"����f��Z�4)u�"b�h]R���`B��W�7~����b_"�fZ�%`��?O#ݛ���S������:��!+��9�N0�)�� 7J����3R뀯 *����J��yL�@22l�E����sX�Y���7B��n}L��>���7I?`-�r�h�����N����ַ���
��7��q�d��!����e{f���N4����ѥ=��֮5�Y�<R�9"<�`�#�Q�XA���C����Nl�� �48������[�Ⱥ��D{�
�hb3��O�~���pZ��.�T�f�*��Kkb���^i9���+�J�*Y)���ߤ'�q�L`���3�sI�n��{ o\��ܟ�4R鈭�uȠGTA|J���k�㛉�QJ�����S/����5����,H��z�_����ʮuY0�D�3�T� ���Z}���}^��c����rz9�熌����L{�	s�酥�Ȁ��0&$����s�o3#g������H���h�6b��BJ�u�<e"���s:����yX�/�j̿Ʌvy.[�SN��Y�����T�8�_ņ�ԇ�<D_� 'H�F��A@�pf&�f`��`�a �:�����,=��%5�6��>p��dWr��p�M���2	
�sE��hv�x�\�?�iՏ�O
胹4X~���<V��(y�:�R��??��4\�Z���p����E�vC	�ȭt��j`dWr��p�����q� Yd���v�У��T�Vh��5ꪐٗ��fǲ<�NI�
�����\F�|���D־`kS�(�uOw�8�M��R[�5Γl	|)���b��׎	��g^���1�����B̰�'Z������t�5����Bi���G�u�)�?[�u�� kρW��u�֌���MyI�<Q_A�U�	�U>���mY���l��,��Dp`GbK$�azm��;Q��؛�*���@5����t�s���jU\��)�I-�F��������{@��hh�WA���x���!���u��R�v��n�?u��ۓ����>� �O`~��ٛ��e8%����A��ے
�)�k�/U�ʦٝT](B�T��X-�ȩ r#`;�/�$ي�S@�B��(���d���MYx(�v�
1��t)k$F�4Uל����-N������(�w�heYbi�.ț���媚��E��Mt-Ԫ��l]=J�b�~�em<�4��T�:)j9�#�d8��B���X�R��}�`^�Wx�Y���N��7z;�Mvq4����:US߭�%�C��0k*�l�7E��3<+�4�'7Zv��ۅ���D]�,	9� �=�%�.Ȉ�
�
 �|���$����Hz{����P����%JK.��o��\LG�U��-0��/�T�� tJ���@��n�x��e�atێ(e�et��" �n�Q�p��"F��37Ϳ�C�y
:���W����i����j��E���/�f��#��ڷ�R�yEz�ٷ<mC�����-@d��C��V�LȼZ����i������Q#������\p��xfȧ���q�;1��3���D/�q�2��g�y��.�Z��W���8}�'B?x2gŢ��h�B���z����� �uOx���z7/&)�x��?�q�.��J����T�0��7 	����v1�V����2 �*���X��2�@���{�_Bl쓚.r&a���ޛݫ�0���fU|����7h�7����6x�u��~�X-*�����Sy��,�p������9`��a�
h��f�[��V���@˕��^�>)���K�i�����3��0���	!�g�)��<FT��KK�1b	qr��r5���9��R�?WZ��@A����6���!�0�L?r����zk�X#���_�%@}yկL/�~y����l2z!��('�ڠ2��ݞ�9G�.LWXş�T�Q7���j�s;e�����.���m �s��=��i��'���o����ρ��CI�k�=� ���#�lG���$�OI�����v��1�Ȑƀz2a)�I���}�n�G�=\�ι� eE�3{��?�|�^e�+e��):)V���^��]�� 5�20e��n��T�8�x�p�;��Y{���������v ���$�F`y.��*���ˁ#2~U��@�P�ֱ����&���`'� ���}���<����r��/��g���Iʲ�Vy����r	`YN&0�W�{NW�v����
����;���̂v�538�st·[�	�<��*� �s�
����v�mI܆�N�n�I�H.��-ݷ�m��օƁ�X|OJ��L� �4���TY�b��m!2�\�>^�[���/e�Cq���E�����r�P!pj)��EPE.{��hk�O6d�~����������Aq}:/����v��l�.�}ⶉa�b�YeI�a�s4:�.���<Xv�gr�L�����8 Ɇ�ԈJH�U��qE�KL�r�1�d��o��R,��[e����!�p}�	;W$�n/�pc�au4�0Qz�G!������s#Fok.�\ߦ�	c=CѢP��8�7><�-�++XyR�L�l�s�{v�ep�\��AxoQ�u�bq��q�V[$m���e���+�@sW�.���C�O,�Of�<T���=N��E�;i���b&I����W3�(IC��?G3�'�/�'�J4l�WTv����3�NB8�SR7����(����>����D�ӭ��2l�P�z�(D�����#��MJ��,��%��׊C�!�-Ka�=�'�<�y�y��GX(�툃��Ge)9C�%�:�f���F���ݖl��F�ҏB=h�nNC���>���sJTbp�rt������x��^t�ߥzZ�a#��s�0���uџ�ci�����W.1���N��Ԟ�գZ�Ko��`E���\�pV��~d�9�)��N�넕E�S����b�.���|&ɩ���q�N�|R�]_�	��RvI��BE�T��@o���*�\x�f�g��h� ��e)1ZD�2��"�Ԓ��a���eQ�W���Y�Y#�hz2V����߂Q�Ԋ[gp�P�rLT�T����"ױݝS$k�d���o���烘O�O>^�G�̇����?����r|ޫ�d��8�n����+Qmr��Ym�P�4��֓��.�]�εv�����&�j~w��BFоt���v❂��V�9L٩з��8��-�C��s�˂,~��`��#�������0)��Pn1œ��ļV������1���$�e�#4�I�BfL�b�?�L9�A�}�-���g��f㯇2^Q�3l$���5 �S*��Y�j����@� LO�Q�g�3�4�{55 O����H`���Q��n��Ē�{ש�>몯meWN�	x��4�)m��%2cr)�r�Y蜇N� N�*�R��c暦c�S2 S�x�%��4�QBW��p�}k'g��W�����$u�H�-��+�X�;Q�|:��ȫ���h���T�lЅ�Y�|}��׹��Kݴ����hs�:��P��=�m����rф�]����|׎m��1�La�r8�_���n����u��G�n�x�Y�������(��1�a��D,�3�m���z�Ӽ�9w����}�s���&�և���xU����W���,d���+Їf_�#��p+���S��~
H?���HG���W�Ɨδϖ���"��ts|�$K�w����Hj��7������h���&����J�'��R���O������<�������e�P�|dY$t�!�Ҥ�������K1����ӱ�VP� ����b��k�je��"���0m.��t�� ��SR�����B[�I�������:_(p�e	�JEx3G�y�
�>̴%���&��$xb��2yX�3'�	�	�3�O#e
��'ti�˪R���ց0�y\p�a������Ƌ��?���Y�rA����F��$0��P7hH�V)��KK�.]-k:S���ARYDI����2���V�Cͧ�!Q,gC��h��i	�eN��z��_<`� ��̷��ͫ�45��?�o��i�ո�(R�ա����b��j3iK<�� 6����0z`% ���m�{�.*��2����˺���z'�3Ns�T��۱�����ʯ�$��	2$H��5����$"�5��`+���A��g���(��]R$Q�����Z����_��z��("Y_�g>Ϳ�2��g(vӿ�^��ڶ�����R�Ye�5贵p�r�y�Qg�Y�[3�?�[B�?	�O�p�_5N2��fkW{g��->;��Kj��
*�(�$�}��ªب�k��?`��v��+O> ]�|I���@!�c5fasD������M�C8�R/� AB�����V������A�Te�+�GJ���!��*ƥh���bq�*�<�j�	*�{�<�����F��y�LS���b�[�
3����:s��F���i�F-͡ `���5p[2��f�}YJ�),� POr?���~(h��7�SѦ���YP@lQS_Ñ���Z+t���ʁ�/L�ii�oo]�O0KT}���g�k�5�Z2���z|͋��ډ�k%x�7<G[�X~�D�1�����1�*��赋���(�V�]A�A�T��e�����B��<����I�!�]|�>H�y�{X�z)�	a�d_��泗��M��Q�J}�x�c�S���Ɣ<kAq����̆F���˂�����b���.[W5�,u�c$UIY3Pzk>�����b@R�A8�d2��i��
�Rӻ��f�!b	��y�Un�y&��S�in��1��e�Nr��c4	aTq����#ɨ'}����c���(�Hl��ix7�f4u)I�ֻ�h��3��X���Iz7+�BJ�ٹv���D�=��c���k��߾ӱ	@ ���E���QE�[��<��%�Ni��{P�_w����eN�;Q��%YX���$�}�xU�7��-o�=a�M��Dcs�4x�};Z��X�E���j�hW��3��E�|)�ȿj���_�j�PN&&X�'hx�_�Ԏ�������>��]�#r�f4ou�*��z�!�Be	�i!Qh�X���F���3�v�"&�-��╡�Ϣ��͑?��`��<tӚ��PX��ٗ�2_�i7U�&�����F���i0���=�l�*0�m!i]��"%��{7��n��E��	�&���ݫ��T{|"�ӆ벼7B߱�#1k�I��Oڃ�!r|�~��<̲.`��ſ��
�1��>�*�/y����RҶ��ǡ%=�g�@�F�_R_����N�V���o6��w�gZ��)�F�����^D��e�c}��υ�YH���/7!H�P�P������6A�}Q�(�5I�o�7ڂQiݯ��ך/�2R#E�kM�q=U�0�2D��E��rɢ��*��U�L '��̐(����]��-\�D����e�ΰ�cE0sd�Rt�_]ckd&�\Pt`^56?�����#����Zd��ZЄ֚��#�w��S�����ڏ�U�y�!1�_	#K������%�k�O�N<}�~��M��\٠+�y2|!XǢ�mae�E%b��FdF��r�
Ě/>�B�u��E����[i^w�0J^�2�᠈��q.yX[R�Z�T1�ͮ�Ñ���J�	���!� pXZ�TL���O���K���N�f�R�,�K0��w㶋�ʁ��c�`�\i�zV�,yM�D�u6���)G��~�
�N\ȭH��f�ͩ�B� 	��FbV3��=a�L�J>T۹�-7P�{�ܳ#��j�W���[����n�����d�l�|*c�l���cv<g�rd( ��]�"I!��hѧ�3��!'�������'hIu8>��=f~��N�>k�?�OG��}�;	1n-��򡾁���l��Nq�K��X�L�-�
tr1�R��`�IgNS/b���͑E��>]�u�� ��	:y�JL����U�5<�_�|DÊm0��E�w| _B��?/R�����c�����8�˷�e��ŋ4�Z�StI��L�Zƌ��:]]�F�l��ge��"�ϱ�w�A|�S�r�SYi`�ԑ&V݃ե�ò��� Zt�F|B }M�������V!r���5�G� /�DH�z�cI�g9f�A�K(m�0xB��:��'tx��1>����,��3��2�ßQ�xc�V��/a�ˤ�qm����[����J�X�-Co;'�ƱȎ*���:���>�&R�=v��X8n���>@Y�9���0<�E�T�6�t�"EM�pLQx6z#��7����kuc��䴳c���Ġ�L�Kh�`��Ƃ����`r�{D�l1l�s���vH,r�TtBeݭ"�Z�\3;{_J�t2�.z����C��8>��\PT*hZF�|FWF�w,?4s?�~+̳W�rZ���M�}g�����i{بXӴ{��׎PN�L��$J����VMP��\���ec\5bv}#�)v�����sn��s���0����Q���fm�U���q�Y�C����E8u�`U� f'lt����_�_��4R4�H��
�/��퀅�CATB�k�_l�S}t�)Uֳ�@�Yz�m���Z5L_�3�Z�~3���p����M�4f�:���m�^�MT��%���Pʛ
��0�OM��.֌֤|rE瘝٣� G��d��Q���0�n^�e��Y�8�x�­m�-~���l��� ͍D������x��;�ޞZĲo">F���R!�鯢#�d��fZ�Oo��Q�����>J6S��Spf�3���n7�^߅Z�+�q�6kF�,�F^�5�,�K�UW3<�L�"�$�$	�>S1T;f��F�(�#Q�!@/�nֺ9�I�I�,���v��}���g&B�-�������̿��5��FI�=!��Lr��W�i}� �I+Y�2�rs�:�z֭]e_og$��=S������6� x8�
�+�&�����@ēcߒ�����AZIf؅����) eu��� ����c��h����RR��!zߝ�i����䁝���k�y�ڒ��-����a:>SL��3fm�����7�No��(h�j�WD��ɗ��i��������>�Z�c*s�2���i�d�[�,�DG;u����V�CK�11[b�>���x�V�Z�-���ܯ1]&����/sqG��z��5�/�֮��߸ϫ{.�(���U�Ǆ��H�\r��;���!w^���I{�(���Ѩ����Q,�a�4`�u�c��<��WnQO��Y-��	cu��{�������RR亩 T�
3W-$�ܧ%��d<�6i(���7A��SѬX^j�鬒"n�ӓ����S�#Z#��n�� �82p^}}qeH�V&�%����@#`ց�z��%��'���u#�`5��b+�`vH��\���a0[�Z��M՝*o�n@�a�G��x��D�S���v�;��9c��`�y��iK.���@�w�>�G&n��\�l_�Ntl�F��˜o)�:P�����w��S��S�*�'Q3��ap�w!S��	�m�N�8;a��NF/��,�.��@H�O�s�2���a��
�����ay��H�4��!�	t�~����Sݭ�N�x����2!�B�Qw�Ew JY�w�"�Se����q�ˣ`=M��͡��_�F'��I �Ҫc�I��'�z�pO�P.�/�h����r00����	����C�Kw40���T��|ͱ���i0�EM���Q�P����%^i��dK%�C�A�/����4��:��<Bw��/���˫�>�0z�ʌ��rEœ��À����0`s������6r��/�!�D��M�t��f�b�����j�1�����XMz�.B��8!;_�O\pu�T���k��2��� ǽ��&����U+��K�3�Ϻ���� �����fA�&�D�~lI��Dz���[�O$�����_�Tj"j�ܮ�taZ������8�g��
��܅.%���g�H����CaJ��-���}Ka����_4�<������p_���	�h_Z/uqmv�N�\H��ͬ��B��5_�ͮ2	����}v9'�2�
���m��D��f*hJ1�y$��frep�#���͂pߋ���4�O5[B�1���e�]�e�2Ҽ/WL��bf)��W��th�� �Ī�'6�o١}V�h�Ib�����S��:����{.�̭T,WI/�y�{,�u�<�l6D
x��p�K[��o'7iC�|��04�C\�^���t�-]YQB�xv�����5�PP��2s�%�y�ϋ�­`���[�R���z�o��L��84{��`������ÕC5��D�yRe����+��\��zFr<���q�S���Z��7�H���t�&c�I +;� =�9̫є�g��D�*Ǳ�-�U�§��nYC��tiL����T�2>��$i���y����`[ s�����9{2[j3g�L��?���2��<�h,�Jb@�3�3ޝ�F�|y�Z��Fǘ"�q��
K�Xm����R2o�ܜpCԐ��6���	jVwY���mϣ@O]bSݷ�Tn�C�3���{۟�+��9V�������*�SA�d��U�P6�P�
R�~��F�d퉖;���u>�P�����X�O�<H\N?IV����k~�X�ҥ��[]?�v��߼����b�Q�>�U�mԮZᨍ������0z���	�i	p!�Q�Z�j��k�&�h=�̄^���_��SBЮ�B���+EOT��Ue@��}Z��ޑ{�����)�|Od�\���O�Сk�B�� MQŏf�z�o�H3��O��ALP&>Y[&+ϾزMU.�/����ٴMπǢ�@�3���s9&�V(���a��u��>ǥ��-,L� ����?�K�{��E����F���\��S�U#8�{��*یT�^������p�e�0�1u��85"��7(��1˱�`g��h��/�E��A}F��1m�����:L�
��I:T���C���D�������.$\[J�k��{�ݷrkO��Usޝ�7OR	��B�[/��`���l���R{a|<��Xy�t�|euc�K�~z1|a��I3! q++V��/	�-#�i�G����� �(����gɥ��^vܐ�3�NϮ@�B����G���8+�d��oS����G15���o��oF�L�-����	��Y=<�G���$���Ca��#�Ԁ��X+��\A������n���ט� %���>����?y��=�P  um��ݒ�bIL(<��Ec �W�3��"�%�bS�"I@��ͤ��끌�H��j�o+���;W�<���V��q�6�QBE�|´}[�\Om�5x�]&B��A'^�Ue��sݤ��<Z����#�;l��	RpE�[�/*/��-�<�\Q��͗�pAɨ��%��ML��3)�P�4�oW[^��U����qq��3�����.a)�~���{�?B�ʭjK�/�lB��,�9�%'�~#L,�P�r|�l�3��-3n��_ <Ȍ>����"R������}!����4�/_�	��Ŧ�D\�&u�x|Z��Ƴ�������W��M�Ct@�@�ڂ�"�ږXً�E��a?�e\��mE�fJ ���9#Oa��f�O����������Lp�]1v�)��ޑZʇuٝ/��z$D��MT�+i���x"#�����Z��bdC)����K��pL�.d�=(y�(����Y�{��������W�q���]>FP���/�w�V1�$��P�twY���ҡv�$/36��>� v�њ��4d�+EJ �]:8��������u��)�.B����[��_�]���� ɯu�m�EMpaL�4��OzP�S�"���fj?�g�2�ޥ�R�W n	�R��ez����R����/�g��3�H�.�O�H�$���&l�/yLz�x���}Q)�oȀ=�*�>��g���>n.`!%���� V���R1�Q����E?�÷�$�q�D�
����m�3�Qs@�:��ܕ6X��KÖ��&���{U6�)n�Q�u��7�$l���S��#J[ !���mb��QPu��Zwµ2�;�H����X4M���/b}�4f�)n2w���%�����{(���A�.I�l{�Zm#�HZ+֟TGa*f����1(}��؀C��sq1��<x�3sH\C������` �����Yj{CLm�E���̨�QOkS��C3��Q���d���s��5V!u�]�-�_rE_�؏i]����+}�����Xo��}�8�,>�������Z������گ����k�1��ቇ�"�ĕ�M'�rzJ2�y�����5h�4�93���5&���ݩ����s7%�D��헄q��tz'=�0p�ik;��S6�Qo� ��+l���E�[�x�DJ�
�2�������e�f��CX�^��:j�+���+$��4���r&���o�Ԝtn��D�9.��`	���p�C�ue3L�m�,�'��c�yH�+F��f�[��M��e�H�]q��KI���wY� K��?9K5�e3n�K���TIXm;���i����B�@gT:�^��t~����G���ʒ�pI�J���
����k�8�0������^xS%W`�d/mK�u �i��i��d�4jՄ,x�_Nf�q��*�$�%�V�,���Dv�q�{�AI��1��./��b;[٪PJ�p�ӷ����
�7�2�MI�T��d�):t��d�Zf;���~�شɧ6,��rZ��N��@�P������P�wws����>��J���:���aٖx9��@�{�ܣ�a�M2%LkT��6�u@<3������iM�3C#�4a_�Lc�8���V�<Y�t>���o�$z�@���	�1,���qj��C~1��?̙	,��m�*�����`����pMg����y��<�����k=�^G�	� DO.�7f��i>�B���v[r�_���g�#w�E��~r� ���0�Z�TfϬeHvM�4g�ܔ
��1ý3�^Q�;��ur�37ǖʺ-  ��w�C�'�����6leŜ������B�WC�u�M8�ṇ.��#�.i�.��d��[��i��s�}±�K�:D��[K�}AwH�Lp����rv����v���I�%"Xo�/3��o>�V�k;������;Z�A�fU5���wi��I�Yi,��;�|�Q�r��y������c���'#cV�7����FB,($���I$�#F�����bYGR����,�p��ƺTZ�&ڵ�!b�s,	|Q� P�Z p����P�஛IN�*��r��>�T.J,�YY�J��gH���e$3�<�TEk���������_���g��A�0y���!�mJ����)2T��mp*$q@a˕`d���VJ(�Ń�Y�FX��f9�dR��y�V+NgK�z�;���� �2��)��������YĞ����+*�UŘ!�_��i��-&��%J��� ���JTw�F�!����ՃGHA����=z�o�0{{�S�5nx�y}0�����5P�#�I5\�b�r����/�;e�I��u����-����sFĺ����ǟH�rE�����`���m�%S�-kk�R�>1�0Eʛ�<��^X�޴f�-�>�L��ٸ�������������\��`p�m��_�͝f�����{g�?��(�������G #2�w���,Ú8F��+�.*�G���Wz6<��:�:z��	SCuڻo䚒ڞ$���I���w�+�A5sZ�ֺۄ����u���N`������'���4���Xt�rlF�K��Ħ�X�6�,��Ū!�<ĩn|�����M��dʴ>	ղX�d"��!�3�yY-�򒁍��{v]�}��t��zU��)��d�p��\̭-*��{����W_�O!��ª��{�v5���G���1���~f�a@�p�u�MW� 5���G�B{.7�`�`�Y���
�E������f�P�d��������=�H�L2��߅*~���W�v��*���fYH�4F�"Z�������n0�G.�Pw �����x͔��F+�EN������O+�{�n�Xɚ��B6pV=�X�t�ܽ��l��J�˽����ƈ�����f�\�@�j�:��'>L�7�������?)�X��L��An��t*ҭ
�S-��HCrO�e�o�L9�)���2�F�OL�j������eR4Mˢ+��U�Uk��x��	���p=QAT����:W� P6S�t�Ue��}1c�[>���b5%Txɻ5$o��|�Y�6S�jS�?��/�s���Mj���yA �$�g��#��B$03X5���\�T���({��&�G7�����m\���_�����$�p񎖥�����_c�q�a�tԷX��N�9(��U��� �J�����K_@�E���u��P�����Z)f]:-!����"��]R8����F��}/�#1|�Y�C��
�$�fH�}� �A`+�:ݥ8��m0�m�� �S/��vV7k�����E\�8��EOs0�L�&��_��{c�J P4c���c�X^���o���CW��s�ka����lVg�/?�%��-Q1�=�+��1�:��acQg��yb���.��{Jr��G��U#���	:��+rF�qKq����y�|x�҄��&UL�{fu��Rk��,:���IgI��2B�x"v>L���6���(:��p�57+��%T~^�7̩�y��|P�O$o8�d�y1R��~Qz���DiQ�ľ��PO�oHH
cI#q�����B���<!1�i��,���P��0D�	C7�,�9��!���^���p�.
 �"��4��?��~����g՜��[����}"�JE�5k
X'���˩1�i��y��*KPo�SFoyk*��\�9
۠�^�Ç"iW-w�->�Z~!���;kr�RHM�T^̹�Y�G��x���q�_g ��&z�.�4��ZJ��W���DCI��Y�EǌC��6̟"'���d0����Ӛ��������fqY�D�伳fW�A�2��_ܞ��U��+� ��i��@�U&��f��[#�?Χ���{�x��qB�@���^fG��A�Z'	!mfC�*�#X�����]���y���̥���#�/������qH3Z�B����i�eig�ȵFR)��Ҝ��f]4[ђ��r+w�q�A��0y���T��˼J�<�o�����{��4���-x�Ac.T%sP)���;P[jg��;;��-�E��A��|��������o�KD� �3\�WR�����d)/�`�T��#q2��ṾL02����{:ջ�q4i��q_�(e��@��3�����2E��F�&G<>�����C�܉y�Rf�uO�$���w\�Cx$��7�B��x���,neS5Nxj9HI)�G��;b� �w����tV�����d�r<���\3j�J:U/Y��q�ͅ�?>��_���Q?�U���� ��A �n�ߍӅ��涜@��&�AY�\D�����ު�u�5�9��t�m,���W�������X�mI=�bY���`$�zi����ܷN"Qyd�<89oJ��pA�>��ݐa^��wex��.���s�XhO0M�|c�sCm��7��H�|��'�� ��(�� ���t�a�f��݅�er��쯌���Vյ�y��5S˷���>BU���f��?T5�N�٦cB�/r:� ���Ԯ�*c|9�D��Z�i���mMuk�T6��.�g׼�Q���	�ޞ[,H���b��ws}ɛe����_F0��������B7�_�򞶕c�}����U���\۸�c`�Ԑ�(���{��'��N�O��N7+O.�"I�wҝ� xlbL�~�l@=(���?�BLU��*p"P˼�ii&"��-@���ˀ@_�_,m�S1^�n�]��TaYH�M6%P��~�\]����Jb��.h̜W��h$pjE
<�Z_���.��Vp5�s�6e�=AVs�#̟��W	
�Y����|��]�F�em92�uA�.v�[.��jFC�攒�Xi_?}�����?�(]E�Eg�����#��C�����e$�K�7bU�yK��U�\o���g��#�ЏfXL���n-�P#��� �f(s`+n~D��=b�х�� 5�U�����@Z�3���f��O*@�)���v�pjuՐ$����w��S���>������F*�E�|:2��~mt�Jk*�w)_t�{J��{���3�71)�z>Bذ��j�±��C�L�&^����~/�����U��>�BO�l�V&	
�������),dN����b�p��I^eU}LId[?���#FaeǺϮ)C���U�U>;�Ü�_�y2Z F��U�ʌ�K}m�!�f{}�,��!-�sB��NH�4� ��i���NN�+fn����iҍCK����� Cg?z���ָ�~�"R{7�o�[�~a
�_9��_�s1Ȋ�42)��W*NE��"M�!�����K4��Ύ�F�r})
�B&h�L�o�hq�~p��}�B	Q֑7w"�l�w�	�K?��������G鹷(�BG���ގe���c	��],�̓���~2w��*��3m<?��:"���^�o��mvkì>K���V��n�\��}�7O�(u�-�����ٿ����ڜU�]��g�b�<:�\R��c��;[�G�M�286'�i�G����:uE���[�Oj`)D���J��H/�$Ԗ�/K��ۙ�H͎55�����l�D��:Sg�5�f���j�&&o���C���=ȑ���d�"�ad�dgMBc�4����fÆ�r'6tS�<#��0~���QwKI���.���$}�^$�	�o2}\RpѨT  �1�Z�{� L�6��
�}�������!l!>E�'��^�0���-�UY�.qxȚ�ڶ�H�f��^��/#_SuS�	T����J���l�c�;]�#�˻�򡺥�~��<�y���hУz�Y��\O�7#��|ͪ�K�	�9\e���8�v�Vw��Q%s��t�8��A��Xx��:Ƭl}E�
���h�������y�]�glF�s>/�=غ��_�V�ɯ2��\��B�H��+B}]�bS:����s�W�}�ɫ+���Y"J�^�\ϯK<h���&�r3�0㶇�J�0j���d���`_9��ė 87��*Ns��xU��`*���^-ŋ�}�3��]��H���9W���D��>h���#sD�k��e�N4�����.�������X�j�����TT؅�X�g��v�ց���b����b�������N�w�v��U*�o �_6��eAִDd��0�ʌ�p��Z��(��yD)�Z4 �yc8��U�f�
p2�p؝ꫝ�/�<�g0i_
ne�_m���G�A~Z'G�u+��'׸r�kk5�J�xg�7���C�b+v�ϐ�ChD����*@L��w�^��l��;�k��P��ɈE��I��F������_��Z��)��QEb�W1�B���o�D�Yi��V5*�V��شp������5�rq�B�ʄu����G�����=;C`4�V��/.�U�����b��+-}s
=�5V鴱z^�;��Q�L�*�X���q:��*9�~k5a	�X�n�Lg�4ڧ$.����>x��n��\�	+�'X�cMM���`�6F�!O��ܧ TA�ٍ����sm��H����a� ��x���?V���m�hsw��e1�W}M-DT��x�H�U�l��T�]Bb2���6:��ڂ���Bf2�|�b�'*'u���V����z�Z~�ESx�8�	O���n����Ċ�A� �;�O�[h�;.C�ٴ����Xx�K�����e��W3!P>]1�0
�p�eP%�� X��.Zܑ��U)�T�g};ʞmVe�C�C3�=���r`HY�Ǻ�6�	��{9&ydL��'�=U7:B{b� Q����?̛�p���m�&m��盨��/���/ڛ�	��7����ۈ i8w�L��}Q$�����6�0"?�@�D��-��'���m��A>�p"p��~�M��m���1�#�gU�T^p�(Ce
8[�.�Z�Ь�[�ؿ?l�{�˪�&�\X��������72�'��kn�c�5��-�#lKŃf[�E�� �]�|LN�\Q&��[�(+�3��f^P��.�n��CG*윗��!�(.Q(:;�mA�8�R����魊L�o0֐�QFX�i{��0)���L�vE���mM�@K��h����7���!:�XtAre�DU=&ߒQ�:�(��H�8�P��ya��ljA�����lp)�/�9#�R?dU�X�.�Yl��i�?x��A�.O�#P��Gj;B�9e��~�w\a��{�I��h\��K�7w	��CV�u���vC�%H)�Tc}��u�Z�K���_읒ؽ��ɧ��ؾ���nŅ��{���,�X��=��T��uH�k-��UX����=do�Ot��!�����Yz�Kj&� �DPZ��Zq��
eA<�hd&���1C3��%:�>/"����H��=/��PLD<;�����h` Y��w�,{���ǽ|q����V��
IZ%!3q8�"��%�;f�9���~� [����w��~�tx�L�d�h�>Pc_|s0iw������F�̹4
>��L�#����n���~���$�q� ���\d��������͐�J�G?/�\�iE��K?с�l`1�	7�c�H����V
ܾ�Y��C��:Y̋���'k��5��B���6��~��� ��C�%�K���GJ,%:�;���SRd���UC��!(J����"��G19��:�����N�=��E}�e�}p�\Nn�ܛ@�����i�C��܁�<*�b���B��ұ���l�R?����7 ,�w�\��,�aߩ��W�5���[	C�Kս8��!} �tc�O��f2��s�[kNuR�h3+�?�R|Z�F�8��W�S��
��q�t+�h��=����%�]�R#2�T���\v�tY�Bާ..P��r���B��05�"�UH��#����BN�|n���hݠ#�%#R���/���G�>�\���7�5�qrh���qj�aNgQ�,"VE2v�(3��A6���)���,>�`�Z���j>�CQ��
�V:dl\,�@�G� ����cE{���p��L��p#���8���/2��K�����L��0G�X�7N ����W��N��ZC��j�����6^3|ɼcK숉�V�i�b"���k��y������I~+I��֞��s�GI�]�H�g�u����E���]{���9�|�M��G5j�'�N���N�yH�n��.d����/%N%�����p��$]�����\��$_�%���ai��UF:VMzPҘ� (��B�a% ݧVu�����U���s&�:�i�����emc�҉b����9N�L�ZR�*�}�,�Q���V*�aP�E)���<�k�@��bqL��?9�H�_\~��c���Y?UT�b�e�ź���g ��,�1�S�A�uu����N�T��9�����Wn͋�be7a�k��@V7Hё'��2՞��('V�dՓt��~5��*-#����NY�H�Ô%Z�`��v�ř�9��$�)�,�����c ~�[�R�2�׾ޔ.��q�:��H���1 �ߖ/�TgԷ�̗kh<yt���Gλ�0"���
�!q��x���mp聣*8�N��{	�ǅ�({l�c7Z�h��W�b�>Y��V��Ն���؄L���#a&'m�g����M�ܑ11z���AD�T��,�v�6|�D�����>W�-^7���z� c����*Wc�m4�L�S��~���]�g��>Y����r�����`<cͻ��k7<�"[�ű��f`8u�<+�y���p��&.��Gʳ����ã�e����m�(�o�/�[� �+u^ߎ�׍�C����˴�� �X��|�����Y���Q~������:�����̡�A��ϖppÎ�����
�<�V�K������}�/KV�����aWC�AW<ׯ>ZҢ�����xy�PtAX���삃cR���P=���lj��Qm�s63�K��M{qk�KD8�v�u>z��y�?Bf�߅w�6�Jz���?7" r��U�GY�邃0Y��-����]�F��̳\�g��Iz�1�
,Ʃ���"?�kB����q�;z� ��`>h��h��yCռ-ܿQg����-A �c�i���~�iR�m�����;"rOU#�N6zQ�6@�:�kx���a�R��A��_2����z ߳�!�&	MB|�xK��/t�q��?뇙�9T�����e�wv�:Up��vhX�t�(�%ބmkÑ�ݾ��C���tAL!�yI�:��K�{uo�� ��9��LM��t�m��~�XA"���ǻ�O�u�z�6��9Pݽ�9}v	��1��"a����{��l��]>=�w��+i�@�'�6��؆x��kw��Z� ����R�[�Gq"��Y]�P�r��.=I�;.SH!��A�5��T0��x��Ě�N��X'���Ы��e��r�!5�-]�t'�ä�S�v_�Џ��t;���1���e:!�T�ΰu	��0�M/��s�̱n5��㙏ɍ_�����ú�S�l��e"��FMT���N�9H<I�jϰ��H����Nˑ�J�a�3�ۯ��?�W�8պ�	r�"_d�j��CD�_6,�Zu��3�D�Y�~��.�7�] �hEL���۹�F�D�c]�\mR�I	�����I�pT%�S�i�b&m6��'K�z)>�\�M�MB�e0$z%�l��/^C�*�o�;��tF������Z�Д�iZG�����ö�>��G�52������k�R或��B�Ɉ��ĳ��������i���zOm�8���Q�h��s�>��eO���u��*a-¤P>|����Jk+�ү$U�x>����B�&i��'Bb1ϵ�Vh'�
�%'�4T�*A`h� �l��%���I6�ec�����y�Q�!��'���A�ҿ�ڭв�0�,���}9�ʝ����+(@�P�7�r��������A�n���3V
���%�mB��*�+��*���5��Db���N:Pa[ �����Ւ�8�3:��ԃk�^���u��=�_�|��#�M���1�8�Z�;���g�C�=]�Câ��/�M�W4"#6����Cz��y���6eI~~��k�bS�G$�]���b-�8tɼ�A�X�ȭ-E���6Ke�K��x;1���T_)7V�s��C��-�����lX�*2��DV��Tr-#���9m��G�[��A�t[��g��lT�hR+�.?�A���bB=3jCk����[?X����q���b��7l�X�+��BO?�A9�]�e��3*t<r��F��χ�T3��]-��t.c����\q���H����tZ^�9���v)��隻g$}sC����u~� p\�h]ӅWJS>D�.�["v齽d-��V�����rc�c�E)2u��׹>B�5of%�4�Fkh$შ�LX<9��D��U�#����A��!"P�q������N�~����IШ,
<��B�4 
~��\2�G��6�ܛ�#KLs�!Q��KQ��t�C���N!(K�nrz�b�0���3=O��M:ۆ'�{�5�Khܦ�|���*��SS����Y�D�F���[.�5r���ր �������: HS�~���E�_Ò��>��$u��������ӑ$�ۯ��i#9��
��V�m:'[a�K%	C���]*���Xߓ8���\I�҇){����`p:���Mi��'ܮ�~I�U�*���z�??�FN8-��FlY	n�,(�=���)���@�)�ږ@���^7�M�DA�L\�`G���)�l��q����z��)�,��0Y苫3�Ps�IZ16������HZ�z;1��п������nI�.<��X��8]��+�?D���+?�C;,vwѭǏ`|��g�R0ӯK�J׈A�=�r���X�ro��U�������r�8�'�h��V�̜�>�zЧ�w>b;],�����}5x��P��ڰl��ѹ���i����>�?�;Z����GS�W�*���Z"^x0f��ɸ/���U�.�h�,M���I)�Ef~w��ը4h8�]T�K�J��%Ud�rtGFBMe���p�|������#�Tx�^Z$q��Ij ���'=�_��}5O�b]��Ҏߘ�]�����m�Cɶ�J�C2�4�Y��Oy�*�:7�)�~���#1�/h,<q��z6Mi��3J�8C4��{8\�� ���:�,Z��Dz�]V��<Ep��*W��z�]50iM������Td����n�g�{���;9#
�hr�X�}!Or,#�y���3��%�R�U_ٓ`�����E{�|,DQ�d_`p2�Q���	��!@��B��/�k�Nο�)�0����M<��44���u`ޞ�b�d�6)�n�eEh:�_2ɿ;��M\� �ը(���h�H�/��=M D�g+�k���H�R��ۿ��v�`�l;���X��s���͸4�_,ȝ�$�i�����r�wv�>�:��N��	W�B�~~PL��0���-wGW˔������M[�?��Z����m�i�)(aF���B������*n4RH~�E{pf1 "�0�'%��s�u�i��\��7Ln�+��T.��y
xz��B@������Y����r�nt%�"������,w�Y�+�}A�f^1y������P�&���"UL�'��rƜ��Y];?�����Q�`��	��Պ8�!Lh���bx�
Ӄ�!'�(}#h���%��r�ő p s�X*�0E���8�+�S���*p��%e7��tF����ԯז�8���A��N�whLL�	$-$��Q"<��~��>@�<
a*���sԞ���ޜg� 2��G� �;64b�>a�C=N���"4�{m�w؀Wц#�n�-��Ȓd+C�7�=2��־�/8c��#,Yq,��y�p���Шc��DJoj����@^
T!6�|��.U�t�^��?�Q�N<����?+�[���{<�4�]�P⺴G��| |迧�	3�����&m��8Z��\�D�١��ݾ�dz�a��H����z��T��:7	���)e-�e�4ڼ�����vd�-P���Ɪȍyg�w9? �}R�Lˮq�JZ����_IǮLa�8+-�Joƈ�׫���ȣ��Ow{�ʹ� $�V��9�c��=��5�Y�1�#��o7�����b�B����Ch�S"O��E��\������R��>����x g&�+g=�ލ����>]g��w� -+����5Q�F�)@OiRF��h��Mc-ks��z��?��&h��Pԥ��!܊-=r�3f�ٚ5��D)J�rC��
��ԿRm(���`-P�n�	*e��]������33
�\6�������V�T���LA�L�e;�%��nXP���o��M`�xc���j����8ګ��L�=^�'[�(XW�#5.�f߶u�QK4�m�@t���iD��枢1�����=6+����9��6S�����z6����@|@��E�Qi��W׃T���#㯾�y̓<@��K�б���gԛ|��[#rQ�8�����e��|иO��ε͡�+3�1�N�
N��x$�W�Y�k��5�hKK�
��+�`��9�R���IpW�.���[�;Q}i&Ʒ���������P��$*ڿ�ۮPʴˣ�N����'���%=�\�m�g�Ç�G�k�����;U�(]N���fZf���'���TL/2����5G�������{���K�)D�5u�@�Q�(l��&||�]9��TsWZ~�{��5UYEZ����}���`.@^-%
1)��	�!"�&����-U��]��;��~�A�i`N�P�a^�%}�͵���>sc�{�f{S�7)C1�m�/n$dLbXĢ�qF�����OD��qN-��8��>4��������b7���VX`(ܧ♕l���@�@j��A��ɬ�H��R{�SH��[l��ޝ�H�-+Gɨ]��z���u�a��ۗ�Ӟ*�م���|!{���$���1��y1�0O\#_�g�E�2)@qO;03޺��fƝ��0
�+���A	�[�5DŬ�l	��IS�K�o�"\( �]5�eq/���:W�?H�����N<��C�M���vZX����9�[��{���D�:����U���I���):�O4���h����dݡ�PO��U]�q������!#nM�F��͊)ޠ��C�l|T���S���E�y�#�	�:e��I1z�=_��rM��rr$��\P��^���"��E���_5��GY�y{\|�}֖)^I���[Ḟ���^���R���Lc�2]�T| R���z� r�>X�p/�F��5�I	Ju��q�)�����G�,���U��]���{v�Wu�k�]�	���&Զ>  �k=hNt���K�s��1���&c�#�,%@�W�� ��E���W��	\��*}"�l�A5OR߼��0E�$'i�l9n��/���������@� �}ԋ7w�L,zpu�
��fޚ"���(;��Ev�侲_��$�[���N�/4ԡx��>�ˈ��}���5�b3�Ev��{��_kC����,����͘E�p>�6�"%m}dx�`�
�r���E%8�Z#�/�a[Ӯ�@��c<O.н���`j�:;����W?��CO�tS{N�o_g*�J�4pԜ���tm���kᄧ��.0n���e���uMc�iu�A'�>�~���˥u�2Ņ�JQ�5ji�X��#�Ui�Gƪ�ѵv������x�R՝��_���F�AIz%���
g&�X~���,�΁������v�(c��R��{�6,mJ��\NG�k����ۛ�$|�m����WN���s�Y�yL��L�����_x"g"!���n���o�o��&9v�λ��Z�M�66'M:���熬G����
����z��{`�-��aH|7֕�v���"G�QX����Ә� oj�ה�H����c�L�1TӺF� ��8�ops�aPl-���͟�G���m��.���Exom���1��JY�)Ў�Y�Z��Xk�؜m�����ig�2^��񡐬�$h�24V3-�nl���Vլm+�|��
�mN<j��IƎ�}���pf�sg�~��,/��3�������u��W��:o������<%R_/� /��z鮷�����ޅNY1S���Q��A8�\o6�����=z�v�;W�ļ���	��<�N1�U�3,�E����� � v"]����M�%�-��H��Ю�.1�2({Ȏ��t�߃��"�y�BH�6g*����aRRA�����fP�x�1h:��R9|H�n'H[��F���3��칓c���\�ΠoQ�I�K�T�I����	C~04.���%��
����C�]|$��=��]��3_����� �wNw�Г�]�T����^~
�#�s�G�̜I�c�����}��2Pe�p+t8&8">�jo��,��Wp�C�o��Uj.���+ܧ/����uD��V%�Z^G����QFsjp�t�YyP���3������-`�xY7�u��r�$�}�JZ��iHL^wOC'H��S?�F����8].Z��J, ��~Z%���qH�ޫG�V哖��\龍�?l�.��g�J)�Y"��r�'=Ƒ,������I��})��<�u��γ��H?x��)�y��W扦�x(k��q	R�9���ً��Fj/�g5v�wal����W$׃�G~*����~�Ց+I��ΈC�KJ�q���B������ק��*e��-:Y¯�^��hY0���ψ��5[�y�gĆT�5� $�-iYy�U�ߥX>UA�����/���������C7��j�p,�����.n\�)Hߘ��<Nu��d�4��˿�Z��H��v����~�]ûP!���<\���1���#j����`6T�VY�3e���e���.Ձ�����{����h��z`|X��}��^����k�����(�VD���9z\��h�hycw�)��m=�*J��3�k�U�V�� "�Z�����ӓP%^9t�8��f�����_P
�n�V���,(A��.mt��nn�#U�æ~_�a�gT){Ĭs�M�!������X*��uLͦ�oqp���}
��Ou]-|JO�a�yd�������ɟL���٩�8Tg?��S��g�q�N�K i4� ��4e��Qc	�S:�*[;]�8���?��Lz��rݞ��FL�G"���t3Ջ���F�߼d��':Y(5��+x=E�Q�	J�&�rq�'/���H�]�t��Ѻ{|G0�� ��Bv��n��43���P45��v=�x�5�$|�UyB�}���f�/yCAk� [V}4R����r�DS�̝G!CK�z���Tǎ
Pj^�J���r�j; �'�ύ��~�ۗ���V���K;ˎ~8׷$�����	��X�m�(ﰰ*9�OG_����z�(�_��-rp��:�$-�BM3-+}�8FL�ο���`����G�B=
�*���:p��8=r���Q�?�`�1�a�~s��su���!���&^e���{-58��e8��QA���/t�kǱ/]u�����J(4�(�|�{�-"e~�CaSBɨ��UՌ�8�F�zq�_�E"�
,+�۶��G�&AW����YOn�����NM9t�k�T����F���/�A�ص�[+�o�w�����p�]���}�C���%逥��xm$�c��&uܐġ��L�+�d�.m�������!�<��)>�n����.}�7(���2,wA��攝�G�v:� ��Қ��_�_k��;�V�/�[R���4�jV��..��|䝡��g�Ћg_߿��sܻb��L����I2��D��#Tb5�n�Ĝ��u@���W�<%��.�Ҵ^�'�X���5,Ѫ}��߱-b��ߟ!��9T�HN{����D<14���h0�Ot�e_�6��C��N�{�ʷ�]�!Ek��Sk��TVƚD���y�}?���68�v7���}p����D%y=I�H+������΁��_����j�?(܍.��Ih֌SѥE�	���U��m�>*�>���=%���펩�3�~=��P�#+)Q�ӆ������Q��QA��N'6YQ�'�a�MJ��M;8kr�b��L8k�<?��	5��2��a� 9+!3q��oKaC���A���������M}xW�����u��m��D	����,n��kKU���J�JL���h`�������SâC�WS���k� ��P[�L��I��Y�� ���-�g��Ղe�޲H�{�J����H�<�Eʽ��>:ڊ��J��fRO��6�#6�9Hy r+*�$eE,�%���"5h�,�B��*Zd��7#�����Ӿ��RޚK��#7+ў�.�y ��b�����2-�2���u�Hl�a�g�xH3W7Q�b�Y���(��e>����ggV�Ü��ጅV�G{#��U^y�wc�<XA�Aq�".��Z���J����׺��X�\��n�"�{�G��c` ����:=�F���4����G�2b�
������R�GO*:�����C��$I}��-�n�+Gwyސ��>�y���2~�B�V�%B��nnz}��~+�I�o�V:�M\�e�_Ec _��w8=�h�kv��8u\���X(�,�����eqC�U��A��Wq}�tL:| ����W��pۇ!!"��5�#���̀�f�L%i��!�%c5-O
oE;�eo��ů�?	�F���O ��F2�(�R�ʚ-�gV��<�hO����ެ�Ezwl��������[�v[݃-z��T��
,{a����D��0���k&��P��q[����r!�P��򁜱&|_�����E	8���UBI�|�j�GЙ����$�v���(�}��)e����
hC�U]�g���P՘>HsGC{��]]Q����[�R���f���T���t��}	�F�F�3�ᝃ�j[���.�;�TK�dek��y`1gXb�k���g>R\<� ��M6����~��hE�)F�i�6�����<��|U�/���X?eq:��/�.L6��y� ���6*�UYA^&ϻk�f߯�ǥxt�ʦ�=R')w�{؇���k��ߏ���d��:��US�s�e�Y����2�:���rr�.�3;��'�Ѽ>��A���(cD�D~n��AS�g���T�W��WRZ���s�l�=��쳎�����Æ�u��#�������7�"�^�B2�zJ��� )�X���Vb#�3����$�y�a�!�ě'����i	�Ξޟ��6�Hna4��h���Y�x�|�w:oEG.~��qbC��F�5>r|�$�x�KW:ȳ��a�)���#n/���ٺx��LU�یA���_mň?����?�(��:�7#�Z5�.R�'���µ�7���>�ka_F8S|�8;��A�=%Ȏ�#8�0��t��J�!R��~������B�B!$��� Q<�֠G�9 �Ͳ���^��҈����s��k�"[3!�ƞw��.��H2b�
�]}A�{���q�[�WrDg֑��`S�Ͽ̾r�1Δ�����g� �̋��pv,y��=�wA"�@�P�}-Rņ�h�F4:�i���l����H(����q�
�Y�d�yB��Ҟ-��,"`��X�q��p2�+��(��jؑ,PT�+�s�V|	�n�f����=��_����v�
x-��&-`�F�>MV��Xb��D�&�X�NU2��\�mL�t+}E�Z>���~��8瓎k���\N��1�Ep@Y��'�Ī�;0��U��wq��v28��"�L7�n��y���1mZ�i>H=�&H��[0u�n�³�V��?�y,t�Q
���v;��)2����C�C��h�aWf�6T(�V��q���>�L$�ȹFp5�Lo�ȓɆǮ��iӖ��Am��`_<t'���#�P?�E��d�l@���AXo�(�d} L;��|Tn�"_�1��0�09'e�吠�q+�q�Y;��֜��v�=AG�ٟ\�:��p�\��X�8y܌�G��Q�_ [��Z�_�13��:��ޠ��y� �w��Q��Og��.�At]wtH��faA�S�z��vؿN�	;)��0��E���wC����t�t��5Q�:9c����&�n�ύ�/�~<$��Yٞ�_��s�����D��IGneO���P�,��=��s�i$w�
�S7t�8����c���FN9���GMc'=�=�B�Y�m��pmXu��W�4W�;����� u�{X��~j���,�h��NG�̣R!x������C{���i�ã}V@d˥U�� ^��f�����גDO͑x��&f5}�r�d1/���$ i��Y-|t�~9R�8��|��(�E�v�sY��̇{���Ode6�w�?��,�4z@���	�G�e!])��|4��͇k�A*��;i���d����2��Њ��/w��� ؑ�XO1�=q��	���.z�B0�F�OT�N�y"=��a�I}Y'm=��0X���X��~�j!�����~0J&+�S����M�r�=+�b��d?���|���|��|ir%��u>v��cR�%��o���C$0U���;�sn��bi��>��JR��*�#�x�^*�� �OH�E�xU���c�y�>x���m�rv��w�/ډv�ySsa��et��zU,/����UnS�OE���dJ)v�-�P�*���z��-�%V�k��`�>$˦�9Z�֎Ir��6�
��gդS�
�O-d�E�v��n2�~�xenv@��ޖ��<B��wB�>�[�i��A��RY����6��uܑo�������^0֋�(TW�Ț�fJ��S�Ln��q��u)"Kay9����+$�6+8�#4�5/ ��g�ȝ���]��#��V|r?�,T�N����S���q���8)0Ӛ2[ݲ�K�cO��I��d�?[����x��������CoÁ<�s*c��q��q$�m���bI��gh�̴��Q���t�0	�q�v������S�����.zt�����%���O
AY����|�R�����"~P\�����g�����|er�HU����p'�Μ3rD��m����}��`�1��_n��ǭZA�j^��KQα� '���.\���m�?�.��m<=5F�Θ�7��~�H��]�92�F���D".�aa<n�E�G�_��@1O�{��X��-�ڝ&9�c\Ԏ�Ѣ�WyN"�9�+���ħh�'�j��%K�;p¦(��^� 5���C2g,��	;7�;����,4��P�&4qQdۢ�c=��u�����Hտg6����#����:�����3����i�*	�	%ynI&P��5��?�(j���]'��u�.�SzIZN���^
E{���d2�_�+p1q.��#A��ϡٜ��X�o�0�V�]D��-��#ܻ`���~�4K�}�-	1G-%5k)$�^ �z!@^�
G�Ց`��������jW#�꣓M�h�&����Rϣ�n4�ҨYy�����j��e�(|:�V ������� y��O�
'�B���O�B~4�����U����=���w͋�|$�!�:�G��[D�Ӣ�v����i���M/ڤ�AAu9^^�r�B��(Uy��ק`�\>`\h�WBSq�5��%��F���
�C�_���hY���׀D�����׸�FA�:�)�n�2D������J����g��x�Z1d�ɉodv��rZ�\�@C�zPb��Յ�cý�*g/n���q.�9�o�S6_���a�B3�z�+�za=|��H��,�U�\��YB�4�و���(���6�Ě�k.�[�7�f�F𼳙_m.M"
�nN���zu��W�4��$Ko 
��$�^�O9�Qr�wgWP+�g)�1\�7���&���9�������� ��H�P �Z�5�0���њ�`���������=b��H-Y2.��R�Ƚ�0y� @��!YSo?�r��ь�"�`�/�6>LGda����꯹�_�GbS8��Z��Q��� ���6U��N��rr)߇��`�e3�ʵ�O�G���E9l�vc���H��\��\Z`��_����L�2��%�4:��������ͨ_�n����]fZ�ͪMS���2��%w�-5>l7ii3T/O�kP�(�Rk������'��Q���(�b���x�أ�H�W������^(��r����<�1F槀�G̬YA�)K�����1���w�UcUg�P�)h�?�6� �=pJB욟�-@����g��_��u_��zV@�ky@C�_V#3P�s��ʐ=�Ghz��iRxق�-?8��
A25M�x��=��J�����*O�x^; ��ԓ�!�HSv>1ߑ�hMX�J J�(�Dy,Nv?xt����G$�-�w�E���7��npG7e�p��)�ֿOJ����N�NwpsKn4���e$�4�H9�9KT�Y��.�Q���Cf$����ɔ��ǂ�b���6�ɵ�?��BI@���qji���\��-���d�s��9�-�����.�pG����@u�_�0_+��+\�/�1I��s͑��l��H�Yg����%�P�F.��	�rg"!�'�@��-�Ug6y���t�$��V=�WK��#�O ��jdB���9bWyN���k��.r䕵Dnp��F�ۑ���q?G�U�����bQ|��Ѿ� (��� '���Z��Pv��|�Ӈ��Q�!���>����r��;�!k�|���Ɍ[ep�Eɕ|�F@�#G�q@ 3-�Й���rH̬m����
r*�[uc��򨯱���(kI�`@5k���������߱pR�X�ܚ�����v6�����<m8[JϘi�M/=��QO`Y�x�Z�X)�O���5q��m8�f6l���0�+G�#�ȯ	+g���5[���UM����d�{�W�YǈN��Ȉh�d�|Y}��_��d��b6���-���+���u��v�s,c(0�%L:Wg��I��(v�����{���7"��N���w��Ltt�zV�Z�(B�n�<�^�l��><�Yq�Ė�u�1.|]�Kp����dB`��K����hH��_x]71�3ȁ��*2h[rf�,�/iL�>g�H��1c�,E6���!��y兏�.F�M;.ta	���&ȸAǜ���P��B7(TEƄlE|Ę�L���&�9��-�H.ry-*�侾��w�F�T �)o=�t�S��n|�Q��p���&��0ʎ��LFH�,(��pK�]��@��  p��p��"n�|s�R�2��/�昬Tc��lE���PU� ��)2ƒ�э�b������{�G�Qn�F�V�n�;DW��*+�����u��ہ�'��[J̈��{�8�nT����,ik�f�Ğ�8��ﾈ������a: h��ۯ��y9_���D�d�S�EO��14*�Ylmt�c6M��-�oU������EBBU�7�|���c������xכ?#�Ǽ7�����<���4�Ӟ���X��n�G����bnŪO^�@,���l���.�E�?�E"%���m��m�j|��n��xYYK��Zˤ�����Ϝ��}�e����7��\�W�/�;�Y���w�gy=Pw��Q]�"^_ʒo��dk0�S�K];Xf��`N[�v���}a��K�q1�mݻiM��6���)��yǴ&d���U�-��d-|^��e�RNi��9qt�QW�������Dz��`G..4Yn�ڳ�j��c�'Z�*�1�e�	�C�q����f ��ql�� �*5�� ;g�Cy�S�{@�rV��Bl(j �SL�Ź9��ȷ�i��������K�lMߜ���n��:�ff����4QE�3�\"�қ�ћ�]O-bH�'�i 4��Y��j~T���T/�A�����d�ެ���-X�b��k{.�re������ q�C�J��=���* ^�nѢ�ag���1pŋK��}�:������ߍ�O�/1�P9Q�����ۣH��c��=�*����6�#g�a}_��7���bU9C|+���q�paߑɏ����^��@��'@�ߐ_ ��l���0��>Ӱ/Ӌ}ӝ읆))��4[�t�	�%fٔ�F��8rR!/�r82�s۱��3�&��M�v�֖�>�A�So(�Lӭ�MI_$����Jɐ>��\��q���c�O���!���6��@s�y2=�a�R>h�/y�b�����v�1����3�1��}� �_	�ܘ)���9d>5FG;N��(>�
��s_�	�d�~�����H7����m7	�}��f��`Z�Q�O�-�V����H�8�N+,3d��ގ�m�z~
���4(���!�,KH��y�ǣ���Kr4p��'���%lX�vZxK[��	�ګ�a0�c�햗���ߜ^�T��f�q�'a~R������*��b]j %��[�YM�N2�~|���t�?�}qΝ�bpμH�ùȉ�@~xǁ�{H�{�;0��8��=�7p���Kx*@� �̢"��$C:���}TD�m���42�{���\�*��}����ʥ����?D�)�N�%���͊f]'Ug's������H/Ti��K�V�3XcU���]�@X��*P��G�4��aX�q|-�D�t�b�{^܁�Z��}J���Gi�����q�A��N���ڢI�4ș��|�`B��L��^"(%yk��ºP4�J��&Z�ĶCt�����'�%X&:�Z��ν��׉�c4�ZD���
ʾ`��V&Q:L�~4�ku�yq�m�D�n�(C�8%�b�묻�K�~.g��v�͐��ty�7�{�R=��2ŋ=v�P��@��?�"�2���?� ��6�խQ�j�O���3�y#m{���Y��vP��g�)��%��>�%K}I��5t��՛ &���J����9 mwK��_��Q�JQ�{��T��?P��Ů�jYoα�v٠�l$̭^��\���;�l
�tĈ�a�=�jJbN��y��j���CHYh�a'Lm9}�z"�y���~{q��$������	4 ΒJ��g3=�$��XJ����d�Ck(8͏���\������X��A��K<�g�]�}��rk��z�#�#���u�1��v�2�ڢ��A��$��Ks��F��~���Z0v�ϭ$�dD���K���ND��h���3?)*c�吡��N�6_\�P:���;��c�zI:Ge`����Df�ly�����2	�L�\�C�~���ݾثU �O����~��@E,ZQ]�	&"[�X��w1Hb;ZZG���,<euq�����JE��$l��\�]�S]�ZNǼm��e�VI��؝�Ky�(oc�|���6>|�@az��*���%M`Є|��cXz�<��޵�A�g(��㠌0Zx��Lb��������bo����؆�3v"��96a���� 8
�)��d:@����W>2oB H�a�դg��(%T�B�C���ǔ	a�;ـ����;��s�� �K���-3�	����jp��&~�ѻ H��o��C��jf�4e��T@�E*�
��Y׉���ȼ6x��q4�b��K����кk�".�e�-��v���E�4����#���Bυ(=�P�f<e������ͭ�l�x�N��+�a\���G���u~l�ZQ&ޚ"c�b�e�e۾dwb�I��h�+l�������e��2Yy���!�^h���,䦔4oKu6]Ft���ERLl>.5@mN.�$�.�X4�(����l��砓|pFzU��*�������������e��\��	�o\���_@v�[w]�`IA.�r����K3�.u��;�8+�e�>$��R:����KA`��8&��h",CV��� ��j,��\�V��#?.��$�CtC�S9�����QD@]�gq�am� ��H|��`/ʻ�����P�C�c�(�b�uI��G19�b�s; +�e�,T�{'пŷeRq���U(;������ZP�׸��j�]!�Qŭ���;4�9?�f�D�[U��Պ�C�D~zę6���j��Z�>϶4AX��S�����ɼ*չ�7�j�F�ӆ�!Kx�ѱ��*<�����<s�$�S���_	KmG0���B�'�*%MrP�����j���h\;OM%��V����4>���>��+�La�X���2vL��r� ��(��hn�=����ę�� d��JBM��s�`���Ȍ!)��fwT����؁�B�lU�*��j�1 ��2���_�3%��>=�!�D�R�`=dV���c�n���� �H�1�mX��M�Q����)Zo�������>�ۖ�-_��n��{�|D���ȄJ*�Zgi��h�J�zȾdM'��^j��f͉����b;�J���m;;!�����y!�u��9C�AYH��1��͵�4�!I�	o����j��{�8̩���mA�sӷuw�x�1��ⵘX��:�~
��	Wt�Ե���ڪ�JV'i�;`��*OCPx4����ǽ73�Օ��8z�>�{�T9db�B�h4���R�d�3�a"�{p����歱zJW`{)Z��xI����:sT�WEL�2�U������9��`��n<!�FEx�E�,.�����@���P\�ۍr�%�j����7�'�9xgZyQ~�4X_d,G�����s�4B��^d�'S��4�A&
�Zz�=y�9�6�����!6��skǢ��2ӱ$��H�=�nNTF��'��a�����9b���ێ7�$�b��ӈ��v�X�W�,��D��Ȥ�!�����+em�&� ��G�U՘e���_-�#8�da�|�O�U�4�XɏɄ%���y��s�{�Q�0�W�ͷ��ˇ���/3��2��I�^�W�`���j����f?�L ����}gD]5�SN���ي���`og��.Ҹh��n�I*a0�)�ȋ�D�m�"ck6j��q7+�8㚽�*�1{�r��[Б~�w���N�H�HD0&�u�%�`��̔�p�"�c�r���uYy���bGo�5���1~���igYz�AP=�kb/`Lh=�� �DW���CSE]|�ҏ4���9J���buCx��oc�۔C��� T�D^Q�8 W�Xu,��=OM���>�S}��|�����Yh�H�#H\��l����x�-
lF����d4��k
���(�E<��l������%dD�j��#v����K�4��F�"j�}�U�~���g�ہ{%��;S��	y��6PhG�]�R)ج�$�Yk��X�a7��� ��U����Ĳ�;�M5n���V kV�Z,��>�]��Yy�:U[����/�B���2�V@S�����GC�t�?қzS�1���0\g_�wS�97�ф���	4�{	!S��tf�wt��x	�~�<KkL��3�e9?PO��Rb��V�s��r�x�N��uǢ_<|YEBd�}�@��o�kԎ�Y�w��O*�Z|��l�üb^)����e�V��4@N���l5�-W���*|?�-�{ ��࿽͞
��<xj}��!-K;UV�B^�����^e�GK"wY��l�������ڼ���B�G��k�d����s�6\q���HM��m�	e�~G�\��ؘUW��y~���/���4Sgޚ�DPy?L�ѷt=��(l��<�9R�遠j��U펥��-��mJKj�� |��(��\E,T�.��6�$i�(�x-jWD�[`�mK�!����`t�����o��ǻ���mDt [��%X]�@H�$�FTB|ҍؕ�^s���D�tG������4�����q�ƝLTe꛻����y�t	4�3���MO{�,�-=��dTlD|�m9K�H3�L��[�Y0^h.������YG�
	��^���
��N��|"U��N*l������u����eg�u_�5�L��L�w�P�v��16�>n�iI����d�[w�^Ƕ�|z�	r�_�����	������9P��� 7s�X�"�D"�A=�Y/1	a�|M�M�uK��j��~k�gB��l���hU�3�M漋���<�H?�'O������?�^a��Z�XJh��;ob��by��O�����1Z��?��}��p�w)v�p bS�Z�{4�SJ�ԫ[�F��x�Ń�F��N��~$·r�z�̤0ޞW@���~����7���'w�{`�)�$d�Laϟ��D�jbV4�����b�a*ƬX���lů�ܮ��O�l�.�C���%����#a+��!ɣ�2� �xm�P�J�9Y�y`9kEWԁ#�����Ne��r�ɣ��'��@<�s��&�K�24;:3�Cv���KJ)���������C���m^�ǃ{y*=��]�u
���I2��W6RD�q�e���-����}���w_@��'�S��E9B��dF#��ӷ�)�g�%؈ �F`������%�c���01��/N��Y��˻�i�����͡����0��jަW��ub�V�5c�Yj�Y��+��<s�EZq..��EC���/���s`�fh�v�'��$X6��/_;$�n/vNK��?��fL�V)���W�H�0�9B�xZղ G6��Ō4�������	�8C��cW|Pic^f����q���3hogV���� �	s�Cn]�ÍAN�FHE8ܧ����9u�cN��l7}�"4k=];��rBf#-V2L�eenR����l�BL�Cu%��P�ߔ���`�����~|U�C�����.�c��-
��խ�d�o�f�q�*ÂWEt�� ��obݐ8��vb��	��@�\��������pK�{'�'�a��/K���9�ԙh�?�T�#���mQu=�lZ�A?��Ni��e�����oF�h�k��Z����Ա1��>�9�#�λ�
7�:����	�$� ����uI+_�6�۫*=�qƋ����K�^�Ҩ�x?/؁sҡ@~E���� �����v���V��ۦ �WL�[3"��bd?���v��W+��YMJ�*��61	][hz
��.�������x���2�޷u��)ӂl�H��f����7i�ޗ"����y�N;r\QwX-��<�X�(+/�A��\���+^r8�h�˵��EH6�����b�aar��Pؾ�lw�5{P�X���o��\��ԣn�^i*�:��lh$�U�S�1�"qV�$w��k���Ri��XRϪ��S���5�=�c\�R%f.�*�xPg�9�(g��LY�C��,���2��x0m�������S�5����2t��Ġ�89w�$�� x=���h����qk~�����rK���4߃
�]� z0��@��Bx�%��4���V�s�z7Y���|݇��T��Z
r��(Fq�Y�a�x���Np�o��v�T�E��+'���{��o�ʾj�(��_F%�3ZJ2}�W��M���{�x�G��o� ��^.>}û�,����r$�0�r��^D�����+���;������W\3$���\{��pp���Aʹ��j�o
9�'q���	�Rd:�$1��I�o��n��1�1��0�������Ô���?�ѯq�3/��s����2
��U�� �E��ݘ�xo43���0[q�u�3��@EG��)qJ(�1�(��@@7��r�⼌Ȩ��!>M"�2ie��	=�B@�m��T�}"2l@k�n�����Mu@����@ ��t�L��+د�����0
�WR�C"�|=`��?P�A�4"����u�wϢ)��Cꒈ�H6�`�7v�]*п��߸a��I�6Bk�T-��d�ھ���Z���s�/юܡ�����/+��� �&�:HjQ�Xt|�gTaQ;n5��*[\Hυ:˅�d!$�j�;ŋilm��~zu�W���'6���j}q��'m�;O�"0٧V�M�Le���yU�EKZ6Χ�=%���%i�A�_/h�����8#̈p�:^
���h`D����}�z�H�P.��Ԕ܉������\�|�����r(��Y��H��&6�F��Bl]�Lc�n$$񢑬u�!�h]�f ���M# ��"��`�`�!��
���淿2��D ��� e-=�N����^iJ�{��P�f �	(KnP��������9p��	GGNBqɝ�R[�-���5DH��q�VŎm-�N���{.�j*e��n\��_�7XNn<�ZL�"'�"V����uCZЙ��8�/:�B����<j�!d�&A�7�y�5�"jˌ���Ia���~�ғ��iW�P��%���ԇ��w��<�	3d��0��˳��7�!隝p�})��+�<��p�:)�-��kϯ�*�4�qT7���a����s��+ m_'�i��k�8�~�"��`�lZ
��%��I�K٪��O�)����M<��D��BL�pGu�{$�+<���M.N۬Ry���V����`o��(e$D��O�!��n���CKF�Y� =�S�kf�*(�'�%�D׬����Q�f��TI �������b	�ډ��E+�����X9���6t:�д�C�Z����F��t���Ѫzo�|�w���/�Oh8)�V�A(&.��`x!��L�7u���6�6^jg��v��o����"/
���?�H�5�b����5[i���b��/�.	H{�U��O�l�|m��z�ٶ9�O\���n�I��x�m��")�N�9��{#o%���Q��  ��Lu�(��	fAi��yHɮ����>�P���s4��cR�_�TT�� ��Wl�'�[L���h-e:��p�8krh ͙�!q���\�e��Y�g�8�iB���ӽm,g�/Jg;��I�0M�)�`�j-zj��,U��AiiqG�hij(����XQ�2��h���e�47.1�#B�d1�tA���g�(K�P���7��}�Ԥa׽�P��'>����GS�(���_i<���y�vPWq�}��ω�|��FP�R��F���em����/vF�w��GC"E���;`��?P%z뼠��w��j"��9G�v��X�Cx2�Pf��.�* 7�3�s^�u/�k?���`֎���a���#��	8�K�1�m ��o!4�}���:��y�H�Q=��[��e��)��(f��?�lK-L�'`�Sl�{�Kܷ��(��q�ؕD���L��F�R�ׂȇۮ9������7����^����P�&���
u� ��.����Ϡ/r N��Z��(ӑ��`��e,��`8�D趧M�e�|����J���X����T�|Q�{�	\��@���8��2T;^�X�L�oTg_�7�����i�]���<q�Z	dX'�+�z @���(�-o�J�b��Y�}���$�.a����)�H�����R5-����b佐���WG��x7pѬ���y����'p��n���G�1^�RDyB�*��,o�n�YJ��	���!�*�JX�غq���|C����f�ý8k�� �cgcRF8V��T�i���"ŭRQ\OJ^�x<0��i�_��ƉB8)�	n��#���PQ�!�e�-q|ܦ����U���K��ߩm��Z��_�3H�ϻ(�26�}�4ȣQ��J���g��W��I:0Y�l&w����(���#��>�N�)�~Q ��q$�̎F~v���[d�nL�srA[L���	�b�y�Gɤz7��xq�&.�#J�\�߱\s:�ZA?�UX�Tך^$�Y�ϗeE2���[P%n#´� �ϓ���H�!'w��0�P�d.28�y��L;�fQ�8͐�z=L�'���x�6�ޱ�d,H�� \�&S���$7K�Xʣ/45Z�J���B^�')NPc��{����汅����l��n��An����%)�;5��'B&zEg�e֯��m?f%#�E�.E���B��:�A��G��`��h�؊&��\�w�Ks��%�jL)�rM�]si	:RI�zd��Ԙ��~��{��BnO����=��`����?`E�����Ve�.��O��;*4�u͈ܥ��20�:�M�p����4b�C����U����[���-���1?�����ٮo@��f�W��3��m�=,�CS��`A���Z/3R�e��?�`��m7���}�Ej60p���! {J�E~Qz� h�^�׵�ӊ����˫��YA$��ط�*NÄ�/1y��;���N��z���9e!��ԜU���&+h%K�+�j?STe`�O&1�A4�U �l=�D�!�I}�O�_;�%��s�YQ�fe"ROA�M���Ԋ2~�pA����*��z�fw�b�^���ô�_S��I��t��I\%p�H�=ӣ��Ɩ�����#Ø6��X��ӯ�/���z�vU�-�����jK�^�|�������&ڷmz�v��0�H�t k�V�[#��馹x'�]V2�2�n�1ep�/w�����\nz6���("�u�qޮE\�R��R6�?�d�Lݵ�wCgD�C錂<WRG�@�����bǍ�) ���"�8ձ�D���X�{XB
o��t�,?O~d"����olm~�x��b��5��@4��hZf}�{���Y�����,�����[��s6��[���<�~�H#᳘�GNqK�	�!n�mL�F|ޮ��\�(��#�ǠbfG~�x�y��7�;2���I��>�Ϭ�Z���'���z�G<�5��Ԃ7�*�ß�
����Q: >���l�Ko2C.�Zʯ��~�0Q1�5��V {���4��n`�9�k6٨~���J��y�R������t���e�W��n���2��)�tݭ�N����x���C���/��g�fz��=���-�T�}�awhN��9�2 ]�
-]�,�/H�5D ���$)����sĆVXa-��G���ON�ұ�J1���j&�ُ�EEW���T�*ۃ�ӮT�hC��}�@�#k�y���Ѽ��J��Z��u6�Ő��5#fE�C�~�l�n4C ʿ�o�_�Le���
=�	_��U���Aޚ2 E2���ik��~���䂴u�sx�~n�4ӽPK�]/��`
��?�^"IR7����9�k�e��|m<��|�2� f���eʹ籵%�~�W"�Y2Ϥm�W���V�iA��뭮��M)��cF L=�Mw�E�1R���x����W�>��Io�yy6��g��l�R&l�
JC18�����Jg��<9�%����ɠ�����CO!������~��6L`�����/���}s�Ql@\1�͊�Ƭ�.P:����i�dqO-N��S��3�-B����]��^3��ڀ��l�-�y�����ʱ�̳��.p(�92�{�L���Ѵ������$O3D��u|�-wP�%V���J�P�#�:W��|��d�R����Uuq�ޱ�Ɵ�39���9��]p�W��߭Q�!1K��9*@h�~��c����Ȳ��F"A����邛 �,i��rU@'��6�<�x�rD�`e�T"�#0@�m�AF��t�j��o�nʠ� ��M�.ի�8e�r+�ښ�K�~�Q�Ҿ�8(E+��KR��kU�c�]�{�E^�V_	���3v�U�
��Hc�_�w�	g�m�*�GN#��Dٔ��Rg�J:��� �U4�-!e���l�']�30���K��e�s!�1m�^uv�A�@8T�s������T#��$?���0�DC����R#ۊ�qB%�Ҍ�"��Is��p�W}*GK�kj;VI�jx�O}�'�
6����P�l�����,��r�;Q��2d��l�v[�$jl_�.ę�bh�i��UC��P�3qeJ�{|�m�k��z��h�U���+u��B�޺�b�0��GF��gԱUu��[UJ���#���,�&�	�>KfT������n!&�"����	ͳٲ��^�b֑�3��$q�$�oX��a�??���������s��">"��G�3�H1 �	K��WqJXOd�	�~�Q�'!���U�c��\��-�Gv��f�����b�3w]E]4[�� l[q�yT�����:ә��ү۾*��쟤j�H��O�$�y&<�;�Hт���k.X<�#� Y�� �v[��&oFV}o�ޕ<4�%a���hc��nl࿗���͌jJ[H�"��v>���ʊϤC����&С�x���b��V4�R�M±�'>/v���G����< t������1�B�oj#z�k��*��X�Q���$-g&��J��C��0��l~�/O��IYO% )�R·U���:�ĚN�?��K�O>Gʺ��,db�	\xm߆�eZ�CUz��GTy/�I��Wlt;G�|�^h}�U��[G������C���c=�0^���B��*�:s�TH��#��G���[-@*uk�:��{A�����SN�R�C!3�5������	$�ࡈ� ^�F�A�i���j���%{�,r�bj��NzC��7BӬw	���:�I��DM:��Y��]h�|�Ӳ=��--?��e7Bo��x�6�'.��z�e?N�N_}q�鱄�Ӟ�����p�(L�+�x�V�֔�K��ڜ��Xz�*�v�d���&y�R6R�O�JERA��(�yDy��
!��no�6�=���|u�F�)>��s���*0�U�����O\��,c���U���'!�m>e#CPV�O���/&����*���PpB��CC)Xb��n+}�S3~R����Rȟ��\t\/���J7���`n�����/	 ��9�O>����
�{1(���k��U�;C���BZ�Ȧ}x��M�'�=�T(R[��
ȑ�[ �g�	�YBs��םËy�<+��g� 8P:|p�Q-��jM����E =ː���DT���P��W��G�����Dv /&�-���hnt6k��m�ab����z|��OU��/QQM��/�_����KK�V����aM���]��o�Zq|c~.l>u�z��V����(ha��� ��,A�]�Ղ�F>gd�:������o���#�qjU%Y^#���{�3A2����TOid��G�/x(C�U{y��Qj����Jfu���l*y{��[�W&�$)#���|x&�v�0e����_����^1ι �)�\��Kvd5v��~1�.��E�Afq0�N'��3J/������1��3��n�kJP;��i��u����ֹ	JDZ��=�t���,��j�✜�!4�oM�N�t���U��NF������[��k2��̢{�iC��	�o^�M�d�I�����, ߨ�4����H�t����s�G;I-(6�����UG��o,L�N/os��n���&�=�j�R;)�_����;V��@�+�萛��tL�@�M�+̞ye��U��	�hD`�<=����C1��_��-�G̺���F���d�`P$i�&]�u�u�%���AL֚^@�G`TzEtW�ɩk���LnH�&�A<ZQj�߰��wXB�	���vї!����(��0��ѹ}r��I#�ϔ?���`�4_Q)�j�OgV�Ś=�����oJìr�S!$x��3o,`WX�;p��SF���}��R���5 ����-���V�uNy�9Ǩ�.�2!��7�,h��ֱ.�+k��{�<�,�s8ʲ�~J�+'�m�g&H�G�Ҿ��`��G�6�!*�E�݀�3x����#�-&�)�iC����u4�۵0�ޱ@V`�A4b62���l�e����+2ST���#oڍ�.�� *�Έ=�j��,o~S����=�,z�l���L��H�C@x�]"�ۂ��卩;�44�\�U�V�يZ�0Do���{��z� ����gDW�
��⸡
�k �H95'L)|G��K^���"���?�{�ݞ�eo=��}&�;�tV���O�E.��o<ǘ�v�U46�mQdֺ�M[�1$w�P����+�H�e!���梙���`���M������(��Y�iҖ������ll�bX� ƽ�mW��&���썮�\t���@�ɇ��t�{�j�fV�^�4M�{^�64.�i�&��@@X��4vG$��OfGۏ0	{�RKfe�8	~��үQ�W d�oc&�<�Pt��W@Z���>�$�dRN��T���k�Z���P�
�ppe�tv(�$���EN�f`�@�2�`l��OA�����$2�8da�@:*ݫ�Q�ì���ѹ�k/UQ��W0uA����ӫ/��PB��Px����E�h԰�V8񖵒����_�[J�܆ɪ��ް	�\�'�.���CF3��5��H,����d4Ӧ���m��i�Fj�;vg�툛K��B�:OiF�B��A�.��,�� Yb��<
��p�ɇ��ÚL�8�����O��~+X��鸢5���f5���ʘu`ɶ��u����@��)�rqʗ��p���qR�Gư��m[��l��]oc��o���fn'r��q]vt�t�Bn&�c���R���9n^Qmm��Y�aY�#)�D��T3qn!�����6���.ϡJ8��&�m�U����LG��H��sZ�V�r��7����a��bk쌭'b'���+be���Gm�~�����+��gp����;fc�GW)ꈋ�*��~�f����2I��ع��66\���WzR��G�bQ<I�7D;�X����k��v+�`�F�i_vɋ�y��1�2�,����*��A!�9E1��e8����z��a�"���d�`L ��e�L��l2��G��\TT��*�ͱK���!dEޝ-��ou�Rh��G���&:	�݈2���qQ��ً�φ���o413u{F�?��W}3��� �f2���n���Ap��Ƒ���"�::y|�-��X�C��K�'��0�=�6�f��nD̝�D��k�
�oz��j������6:�bԧ��� ���GhV���Q��U�-��SX��h� L�Î%����5��.]XkYO��r�#sӗ>쑲�����Ǎ�Y$����e�ƬqtH�$L�)����ɼ�Ю�~�3c[^�q�I�
5[@��ʴ�.��{�Y7D;T�Pf�kj�8�B~ض�]YL�G��@x��V���^r��l�Kw|�#q��a�5�f��O��F6 d̪�8��M��ð�C�	���[�*�f���2]�~�.�8y�$D>�� �C-�������'�W,�3T�B���oð��u���1��\j����}�<��m�Z����º���'��P^���
�K#���Մq��b�Qk�3�h3>r����@8_��k����L����?�é�� �V�oR8�N�/��V�������$��t��+e��=r��͊
��}����2X|�OK l�O�B&�rp���Vs�1��ש�U����:n�&��C[��ծ��Y���a�z<nLZ�l�-65��܄� Q�����}e���I����;����tC1>U_�����Fk"D&$��4����
�1P=k:���ʨ�J'��ok� ���t�|��z�i���ل�sVݶ��F����:r^��*�r�Uz��1��q���`Lr��������U~Z�~_�_�v�(r�~��r��Zz ��}��ue�u]�FH�SX�l�#�2��G6����$�����r��I I?{4���myEԿ��@���1AjD�z�y�g��E)����,�m6��*�M�aInUrY\���33�\(�"5e��{�Kr���2�$��ao�����u%�*)�7 �0�z�����*���xC�)�|]�iI���jCW�_4�t�D2�~េ��;���U�R�������p���w>�e>�������m҈�h�+X=���=��A'(*�1���~8O��<�r��D��x\al���蘶�\ߥ�[vNC��}�{h��u��Md��Щ]pG���O�����K��g���7���S�aI��[�A����;x?E/.��Nd=�R�mM��5ED��vFS`�*��݌n�j�I�����z�c�JsG#N�$m�W�<�6�>�N�ќ���GbT֝���֝��|Ҳ�0v���ؐ���c�m�%�$���iv�_I{1@'Z�6>T���9�c����b�h�/���.'F�(&�JO���;��؛�A{i$:��ds-�J�BQ&^��v�vy���l�������>+&��;�-�b.���lo�p�����>��v �$ԟ�7�cC����F'M&td�TM���P��qD���j\��҆��.��<�p� z��MV��Fs�w�.N���!"}�U�x�'
ũ&���p�����E�G;���1r�WH�!ɱ���t���?�{�R��늦g$�@玠�vu�à�ѐ�5�㿮��H�[woN��]����yy=߹xn��vz����~�ȹ�� ���3�h_���Է	#R�.��
S�	�	��sT!��6�a��tc5ȑ��\�;SRZ�י6B�i�(�@�0����=(#�k�h�a���!?oK3�q���f����P����¤=}�==�9"�|Yաt�W(�=��B
�_��&�-���X�m�>��:#�}��Ns��y�$�Z^�����_�|���?\�|��~n��H�3��ٍB���OzU�����)$�B#���؇�'�db���z��Ap�*&#+��ɉ���B>B\y��x�i|x|�'||����E����%CV��{��$F�Z.��~�x��K�(���"�z��W��ԛ �(W�x�M.}��5���yŹ�@%�`�'�n	��Z�Iq`i�c�|e�(�p�%�f�(��,���ˆ���_����,�|v�OxF����Դ�ͩ|�Y��L|}�����x� ���*��9��C��� ׫]y0�ҕH�G��S-\�Y�\U{��3�n䢿{�R|&g���a�yn��V����@J+��/a�*\(B*��fT��}>Rǈ-�f>�i�$�k��p/�=��&fKX�*GM�z�i걺^Pi�����C�Ve�q����6%�/dKe�I����uklJ^���>�yO� �v[������:l������w
�#Q�Y�	Y�<x�ѱ�Z^���s�!ip���wo�1�s��N�wp��;�
��g㵮�_o�^�����C 6X�U�gȫ���T���<�Ŋ�"ں�W�q��e��G��DE|�S��Be�$E�x�s3��1��5x`�0�UP��_Б��/��2+�:�f��N9y�s6�_v��`0-���H�^�W-����Ĭ5
��K�!�g�ڤ��ݛyw����&�y3��P�~��T�J��m���Q��Vx���\(	P��<�&�ُ-�]��)`�0��i�9W����V����\!�_�$�����y�@,����s��R�@��nl	����~�0���eSk�s�_��_wi�H�20b߳��cC�� �Z�pk�Q�'/���a�!���y���ߎBI���:���ZD���������������DL�MH����)��8�!g�'����8yZ؎�$�1�6� �a�����5+���jHR�e!���K=&>�|%2�w���Z�ԫ뵟H�l��M�m�}֝����_�F��C
�+��(6���(��K纜c�aZxl=^��W��W0g���?�q-�A���n��4���7��y>n_�-��u��T�i��ő��N��[��G�K���eJ:s�|�[>���c��m�u7�b��iNl��/��}^[C[�E�_]��w�ڡ�tU�ӦĦ?����:	���W��ZI�*8�*%�i�?QU�ˇ��u-(>h�e� 287�2!�+b�u��~��p�;5ƙD��r��2_��Fjqw��{������t,c�ߺ�����>�V�����͈���^��d��`у�kQ;%�'��0<��GZH{�wS� 	�q�XM�/'f��[{Zc��2�����g�o׈�3p��^����A����6t/�⍅���x���_�\$�s&Y�봬췻=���ɘh�3Gvd��� 	�/ a�-j"S�w�IL�ui�,���~�Y���֓���2�]�瓁�Ɔ�uc���7�佱�<H?�����3�i�A��$>i6ׄ����aK�T&�"ZA��Hw�n�Q%N� �/��x�Lm���{��M\��Q���K9K��
�$~��XO��є'�MW\ݐ�C������Ȁ��GF�����Q����Bk�T�ٹc�v���7���2����l������������w8�O�+�GH ~��+�L~�%�T���W��PFz��f};��|[_#j�j�y����@��F��J�rQ�S�HHUt��2\>���J��{1�=�*�q��H� �1=U�E����Y���M��B���Ċ`�����j�IyA���s���ay(��GW:�9���]�yG�In�n[�ɶG"'��8$(��JANm�o�߸�v���Lf����535���]/��H��	�[ ��R����� 0��<�|�y,/��g9�����꫽=̾�d�kyb_BoyvS�/�QJ%�Z�u��c����f�r)�i�^׳�ޓDIN$���ߊ�����G�ŀ	�"�|�W%l�P���Ex�p�q^D��B�!�����N�$	��Ђ�Ԏґ����t�&p������d�\~�'5�Q��ϼk~���n�#|����I/$W�:��] OC�a�r��O�;��`?�{->DMŶK�-�	�NΣ.�������E���!i�I���gU�f�����N��Aջ���0x�,)�|GF�	��$9f��ZÁҶB�?��2��L�W0:91J�E�X��w�j^�0]�OՋf6T���D؅�1�_lw�h˹l�j�6G�!pX��w��0��!/�v����SE��W�D�p��\�U��ra [zj�Ncq���*e�P��H�z__�z
������x�E�sY\�6$�w�@��j�^%K���c����Q��T��m��}���u0���j�`I� ��R1û=�g�֧n5�&��c?�H�<e�.�;t��-uecj&��r�ek�����A*s9��q	��%�ED�/*��/3�UT�`��{�FXX���vu��Q|���g����eE�R-�� ��1���c'��V�|�]ԔYeW��	M�pM�co��\yb?�3����"4�ɾ
'�a�/�X��В��wW(^����G}t���F�Bfi��Q_,��)%࿶~ ���H�\��A�b���@��'�v�z�7��g����<K��ñt�zge���ܯ�or*�jL"�ջ���45�/Em�ёZ#���j.Ι�V�����wF:�A����n�#5@�>\��M\���!��<��q��g��Ҭ���Z���@��5pi��M*�X�W�Q%r�G7a�b߬���xV\D.ܚ����Tq�+Io+bg�(�C�V�$;J��=Sި�/|uw�q�%��x��qY�*��VI�ԇB�=	��i!��عK3�*%LF��~e�?��^R���]ez"��Tm�]��Yw�V�/����t��ܭk���L1L��ǔ�^fo�^N������r����qsQb-KiW��s���ߎ�(Ç��!؛�#����N�ūɞ�ǒ��hw{x�*�:��z$��<1k^�ܭ�䘫2��� ��D�gK9�8OQ%%���a:}�0��"`�d&i����t��'Q�`҇�����V�ԡ+���"�t�,��6J$.�����p�E�+�!��5��BoRFr��#��~8f!
f����dc��|�h>e�\(�b�T��$�hF^[:�Z�1��%?tu�t0�@��gTV9�+8����������;#F�a71Qea���e��a:J<9�D7A��bDƔ�Kg�Q׭��"����a�xꎾ�[����R�pI��3-�������&#G����L��������Do�s�aЈʤ��	����
��㼗��~�}4:��?u�θ�jR�c������܍{��!�7r��U�_� ���o��]l�SsB�8�P�^��0
����(�o���|�Su� ῞��U�d8S�rc�r���nŶM3�&�D�y�B��B�G�wu�>�����xb���T�v $�r��AdZ��N�t�>wq{�������=���M����'5
�o|���`�Ё/�
.a�E+nkjz:��뗫.�	�(?����P��Bh�9h&�?v�z�nC��-@�2B�Nz�0����=�ʯj2G&ʠ�Cem&+xgo����K����w����4���>�r���hNlom�z�@�w�&O�����Z�^�����E�)������� a�H�-��}8���@#>cT����&c$_�:��37_��k�������g~�;��QQ&Yn]��R���U'm� ���a�E�7}����!*�"�i4�0�C%"�5?F��̴�U$g��j�/�=�����O�3�Վ�G���?��;��p7�$�w���0��6)mV�d��4����.]d�����n��Ơ1,���B(��k����DZ�:ڛ^������R�Z-LNh���O�
���1/TD8;��1���EA>D��������R9=钭`�����T颷>H�c�(G�pX���^���\2Q(���Q�Ӹ%o_�ϩ9x$,���:��LV��EOh30����8����Z5��-L�<m	�^4���yq�6�F�YJ3^C���F�za��SW\�`��,C��~
��*�=[��}��pJ8�q��M�"'�z|_.W��3���)2j#_�W!����`jE8�y;[{�ഌ�_�),I�s�щ��s��r򶷰�Y��+����]��+x*��"���Xerּ����w���	�����'��ɸG�w��A>�=��B��d�|�䶔�5������<���Z}6��Y�"�\��	���wi�_�!-ow8��~>R�hj�J���[̬�:Y�d���d�G�<�mN�anu%�,ix�D��C�9<k����S���S!�N�oR
7�`��k�t�C����(H�@j�W�[}�i�W)�&�g}9�Jˣ� I��&|]6)/�x�?�x'����[Ypp(��W�Q��_f�}�Ľx�o��4��v�#5��I9�'L��@Eh�Oӳ������"�y�ݾ4?_g�	g|�-�cwO�������~�� �&�?�f��4.D\��*�vu*�X�Y��Ղ��ߘɨ�n5�
�r^�xW���-�D�'94������
����2�'�ы\0R��UE�Bp���og*���P�0vFl�9�[���DIEPƅw�!�:+��
С���w�isN�[
�ɐHv wB �H��d�Z�E��s�QB;z��~��
�x*�9d��z�>7��M�'�)G�vNOګrT-�!yIcyڳ݌
9y����G�X�;��t��QۛD��������!''��_�N;K/�;O-�vK�@p��i���x盅���y�8Q5���A�e�Cx��>c��GeL������`폡���m]x7��:��Jݑ_��\�<&@�������C�r���-�#o�7.L�c����d��b ��>>��= �R�Y(�/`�qr���f�'��!S���h�c��o銇�����o\V沸�8�9<�g�wS��;c��6��J_�� �g�Z�N�h��I��5�n9�S��Y�In<��D�s�c"���ڝ푦s�&T��[����%'uEW˅ogD��'���s��4��w 4\xP^�	;�xjYF�<�N❍�|ĸ�)��L�c�֣]~�z���[�['�T�<$�'�u���鍰�)�@�v�Mjd��	�7�s�nHz�8&�W����<���r`'��|���Eў��sWk�yzPr�1ݿ�)����h/��GS�Q+��,�L�y���/�6�x*�'��Vn��
<-�^�k�lៃ�|����A",��d�b��=Z��������2-��EP!ɕ/U9ѫĽ�=Y,�u3,���0+����ڥ������&e����d���E,����Ѧ^��p��^�Mc�1ƃ]v��܌2�N�{��7�@ "���t���xt�<L�R�[;R�N��!��\^]�Q�7�U!�T��K�{ےҦWs��0SR<���&��y"�K���;ᆋ"��pMm���\�=�~����C�ٷ(O���>>fp�7�`m�]hԲ���rD0�"��k��g�1u��})9�ڴ�0=��l^�T?y�4��:&X
$O*�w�q���8��a]2M��2?k���6�}\��O �I|�Pn�����J] �Ӫ��~<S�����r�GݰKu���Il��l��.g��N�y�^{Yl��`d7N^M�����,~��c�{rHB��.Ik���th��Z�k�7*��x�a���.�_����ۑq��UWhq�_�V�wZ�+V;�/���w8�:�v���E���at6J>��9�<���٨%$L\����M+�͚�vf�m�gs�t��l�c��5�Sr?��:v=�}F���G U�h�\�˩δ냃I��I��<h~��o�ԩ�Ek+�\8u���W;NG|Y)�2N���7rMqwؔ?�n�ԅL�E�O���t�nXiK��C`�9͡M�qN�y�"��zp#ӿ�8T��F��.{~�o���;��Jb'��ga�_;|�e�·�;"��~����(-+�<�׷.`{Y�%?��Y�q�w�c/�6���=H�I*�۳�`'�	��?Fb3�<85��3�z����q���e#1��	�����A�<�#�Z}��GV�7滖����Q�b�y���M)���'*"�6��C �RQqO�f���<�����;jK��f/d�b�ŕ{{ԟ�aZ1*,P��~�޽W�0{i&h�rS���tDCO�����wD��<��
f������B�"B0�nn�8$���ݔ��F ���݌ſ@�H��8Rk_��neD�Ǖ����w�M}(���p�R�[���[l3?P�O� sw&,@��D����!.ن�9s�sjWW�`y�Z,���ڧ�gZ.�-2�"�����I1 �M�m�?n�s����!�;�kg���<��,������H8�qw��|>�Z��� !�6W�7�������_`ѿ	oJT'��&ba�3�:�l�pĶUt/}�%���7<Kir6��8$GTs#U�qR�߹�<��)$VTN������f�l&�(Z����b1Q�+�sf�����C��a��˳1�G2}G���o�oPϿ0����y��c6y���ɤ�1k;�%���l�TÍ5l��E
��_���I}��9YZBi�U�X��9��0le?S�[�� ��[�6��K*	������Q$���(�[_�hN�Z�*W�S�6�����=�;��;�����҈$��Gn���>֤+�\L�ζ�3��áΈq��+� MT[��������P�2-V�	�_<�z8t���{�#�'��Q/l���Jy�V��JK�U8������u*�(L�_ۆ��/Z"��-�5d˞C�59���>��몈���j��*�L�����1i�_��3?�l0�:�t���h̻��+��.�0j�Y�{*���h%߮?�8�!�{�-P��aO�V���~b������{���E����A��8�<˓B�˫��f׬�FM�"ְ:��߮kŦq,���Z���R:xx��:d>�S�N�����'��b�����������yA���Ӽ6�3W
��Vw��=�9x!�m���&m9�>���N�c�(>dr��Էû�,�}G�O%��]����;��TӶ��'�W��E�N
�:��'i�I%~�����M�%0k�[�V�(��o��d\�{���Ɛ����ʖZ�m�B뱠JG����j��-�(R�4��vÍ>y�{U����(�n�xT��4�;�+��h܎�ʥ��DM`���ϭ��U�hs	�+)�)�Vj���ۡ��p��K>�����^	��2����Ҳ�� f�Eu}2N�6����S&�N1�m��G�l��%y�xx�����j���IPONw���Ț��Y���w@�/������!�v�O�PV'��]��8�tԓ4��4�,p(�Y�f��o8vpy�H#q�H,��F̭hXv��c���Y��Ky�����HSۥ�6��S;����sT�������S�#w���c.v@�B��I��߹�ɍ�G�g���ެ����+���{/������S1��x����@�>�G�؋�b�l�m��ի�K:Y��H��<��u1~�3e�����9�s�OPX�^6D2˽-D�zҋ�W�2�P��ˁ�3��BzC�s��١ʀ�,j檂 7W�B�lQJ���� ��/���z{�0H8r{�ͪ�?���D��m|�1�x�g6�K�ĕ��3?�@IaOm����)}O7E�m6�_�eH.�u�ξ��@�w���2��'# ��$8'2&��n[�p
d�F3w��2�Ƭ��C'bS�w�k�Oi����)���>�M�O.w1R����AO+Z��'�BK's���i6ǀ�ƙ�И��S/�M?�0l����Ѽh
|F}R݋ "G���,ɛ�^�SV��d�p��.��|O�l*V�~2J2A�24tiHo�hl��g�mܑ��揽�2z<�3 ��^M�>؞V4s�V�ײh�^r�]R��q�=nr�����[Ch�Ze9������DB�л�/�9e��d5W9���z�e��8��s������턐�o��|yM��,72���
x�R����{	�Ut��e6�RH#œrt���Ӷ��@]�%��R��u�W��#B�	������:��pbT��P@2?'	��W��oԃ#���8\#Ψz�^>>��rqـ�.?�qH�ӛ���e���IMQh�D�?"�:uʧ�]�,�bk�&�r���Ўbk��ۤ��O��cU�|�#�1��<�Q�z��n��r����"��7knK�jS��p�ߵ�j�;b�+���f��$���|\���'��=���������t��:��}����@�����g	�/�Ţf�%YW�]3���j�ҍK5<�Ԁ"$^iz#�ܞ`�c�F����p�
����rTPg��7�ebņ����,pS�ϭ
{Wq3��
I�����Il�
���J�=˖G��\�4?�_�##M��첏�k�\�t���6"����K���KJ�"�<��hI�G,z�a��������X�H��N���k�9�Vl-��`a���ԫ����`��8��X^�����3�+>P�4�z�s��T~u���\c�dj��f�	��(|N�݉���9�q;��ɉ����v�����I�����(`3&y據�ecԯP�F!�Wg��'�a��UA����)�_�̞m���zQ*{�v��ǭ��&��B+�!�:��a՝e��F���$./�ɘ�hJD�������9�"fNW��*ZDlW��t(�]� Htm/{���Z�$�Q<�o±�,~�L��O��w�Fv4'�"3Ə6�K<R�t;�?
�	��/k�FS��������6���;Phi�r�ۨ��m�{ԅ:�@�U��GV��:;z�����n��*��=L|m�ԏSqqH��z�m%lqr�M9C"�n�>�������l`�Ս�&d	ByEԀ��B���1F� ��ٌ甠My�q
�J���x;_^t 9��K�8@������P
��O��3g�$��ԪV@�
a��>D�5O	-ѳ�HbW���3.>r�������4�x�o� �x�H��Y[y'U�RO4�V���q� ��5�ഞ�<�7 z�6'޺;��b�.��9�e$�1.Α)K�-&�K�.#VK���"\�/IF��S��"i�!#����3Z����':�Vۮ�!%G���"D���lI(J�E4������qZö�'�Y������JP�l����*����͗���˝wf< 6q�T2����Ѯn�0�L@���B3ʶr��J�Xڽ���KH~~�!E{좿L
�(;w":Ώ�/��W�Q_� ���2�F��&������Ɉ���������~a���	�k.��yb��a�	���Vќ�+���$l�wdM�z�ѹ�z�ku���Q~����r���j�TǺ���	��ρ �wD2m�J>��5�����UՖ�v����S+(�'��Z�:�Zߞ����0d����u��,Ub/�;HT�X}���P%qG!QR�R��KV�BپP��d�]��d�R��U���� �����hUg��E� �H����j���7yk�R
����z�'e����ş�M%��@�����MZ�hzqc�����Dcr/�����v�C�&M��D?���Z����,y��c�	wT�e}8���]�s��4 G�j�f
^`�5j��\��P7d6��x3e��t{Ta�Y2�+�&=�MƗ���R�c��}ʹH��.)�>+��F��ġ��4�5fC�*�%�ࡐ�"����lUsO��^��S',�~'7""Q�3�Æ�(Y��\�t�|����п�̅�2D�7�0�j&��š_p	k��{��(��A�7�!r5���I�G��ȩ�D��GW���C��m�{|ן�"ùs^XQ'W��-�jR�=�Lf`�**��LEٹq���<�0��Y]�{;� �+��~������p)]���Z��+��	�Ȅ�Y�L���uw��} �=�3J��i���_�Y�-r��[�x�<�~�jB���<쌿:�A~�
!!8]z�x<u����Z�i�O�����,�	���NYR���ĴQg�E�0���ӚF������"L9�JMHC��* ���d��z���ױ*[^^k��U��ߢ��-Bf�K������
W��R^��eX �yn4�῏y�#��;�ډ+ �O<��m�wD�}Hz"S�"���K������خ�H���/���%�$}��� �4�'_�������B�^R���XbG폂#���J��w��㾪��#��:����N"�?L�Wz 7K�/5���1�aB�A�.]s�4C��ү+��o�p�@�o��啫X�;2�9�(�0�1�,5��m����QYn��^��J,'9�����T����.rd�W��7ˊ䝃W����H�
��9$ j���v��W�H"���ipR���_I���2����9I9e�l�6�C݉�d@��u讔U�3+{����W�^(nIܣ�[3	���͊A]��vc+�R�YՆշ��QaM�޼�g�z!}"hI@�/�� ���d�HO�7�w񍌠��^��!u��\�a��UMQ}.Wb@�����R�$g�W[Y�$9"�l+ߴJ��^�������r~�v�ʀv��iƗ��oU��K�X��x�a���O��$�YÎ��蓋�����+�5��V2�1�2��gtǐ�<������h�^k����(�ɶ1�W���vw�@Y��n��g���?�q&%���_�c~�L�^�r�2�̺�~�<���-^�\rE��>�`�n�w| CA���
��t=�Pӷh>�Ǘ��6)ˣ�b���E_�6�"z��a.��� �O����t��)n��0UΒ�!*�᷏e	��kA4�P:�@�,`��ӧ����Ə�V����kP�ｏ���f���D�dR�����i��Ӏ�ᴍkܜ�j�����wWؤ�����K�,�6v�<ZL��e&��$%��Tkɹ����j����y)�[�G��o~j�J�8���n�����Y��2�i��k�:�@�5��b '��i��?2eqd��^�8��r&R-�B�s��t�Pۂ�5��F\T��cve�1�oV���sْʺ|C�>Z?��y�ߡ��P爂� 9V�)�C�y-�;i[�{��Me3�����гm�HM��h�<x���ހ����u��ytBf�8�\��ٕ�@�C�zAM=!-(IFQ.��l;��3;�Y�[����:w�l�(xH�4U����A�w�AA�p�u3 �n���;0�دE/���qq!X�� <���T��Ws
�e�I^�E�?/�j�ЗgzS��^Z>}cG��Q����5��ں�;b�7+���IXXp*`�#�H�td��N=`�H��k
>��#6uTb-�s��I�vX��`�h;-W�/����U	��$�"��7��n��@$����ej*�i�i����n�C�eBvo~!��m/?	�taU�����2��v!��^����U������q�*�D�h�wAR
y���4K�M��ԥ���#���XE������dv"DnG�nw�g�|�t3μ���O\��~��7�0Ӭ�T�85�*�>�}M�
��Aiߑjv�
yM��z�Nt��
���|�^��k㲼��+>X[<�$�%�K'�̬)�5� ɳ� ��/wKCl�:Pبj�����Sjk���q�$��ߞ+5�$��)�9����UrZ��<��4 w�,�E��|� w�yX��ָ���b�D��id��U���9���.�D��逪��W�R��~�����$���U��z����7-&�h��$�_y�g��@f�����e��e��j\j:ۮW�錁��"m~ݍ�P��6�Ľ���2������Z�y�f�WM����.��A�M�~�튉�c�͞�W��Tr��jc&$aM��"S
���8WU6y{����p��0�/��z%XIQ�$�2Ń��Orp�il�X7',�JV>�[�xҴΪҵ�CzQe澫�a��v�}J��=�^~@^߆�$w*�	��O��`*��;��1��ˏHse��|f��ib�d倣�'ج���}c��$z��V�ň�[��y\�r����HC����-����A�����g���f�T���҇�f]��X��<��p.�
n�����$g��^�I�u���?�Z\�?@0�4\�5�-a� ���9D�¦��O�7hU��c��Ҝ,a�HP ���`����Y���j�7��_:�*�]�nW`n�PۍUX���s��n��E�SΌ/զ���w��VƊ5�.{��Zl��30��%՗T��c|���O�_Zrr-�N�s"o�i�B>��bs|�����1���K���3_D�q����z�I�<IЎ�5�v.4�� �ڨ᳽��B��R!���������[���hh����E~��ݝuE4�Iz�-��1�MXMDr)�\�i�.K �G[���jl���*9�.��-	��ϤS_8s����Wͺ�Cb��ᩓ�$�~�ˌ<J"�KL��P%Sgs1��$*���a��%���?���a|7[���[2��}]u����_�`�1� @)��~#{}��D��@�yS�<�����.�����L���[�}*\�S\_Ŀ|W�՚$�+�����[�Z���ʅ��ö��YU�w�}S��v���F蹳	]A�5
ѥ!��D��?�P"���*t���e!f=آ�mtz:��j��	mʤ��� �%���(��R\�k�ka�?�`�D�h��O#`��EZ:P�X�w�����R;���D�aG7Y�k/�s��O���#��H4V��=���FA�_b���x�͒�(�a���"��&y.�dO���wR�xÒ\��"���u�&�kӅpS��Q$ɢ��0$tWs�Mx������.xQ���R�M��[F]:��_�S���G'�	7JU(�h�����9F%F"�V�9�e*�������:�5�TB#���0u�2i�D]�cm+?�c-E:B��vF��A��$��[Ϲf&��}�:*<�U:��Y+�e��5}� ��Ԉ)f��>k��R��A�oޘ$�U����LS���gY��f���n3d�ևNb�E&) ^TD�9��p��'yA����)�����*�FD�e���Q��=,̜0Bu#�p 2�X~��?h�̧���ca���#)�+�M��$�p���{�˘�#��X�hJ��.�[����Q1���a��4| b�[����L��ˉL.�=��'�OCg�r��I�T%����`�z�����1���LLm��(���)���̢ŴL٘������2�#2O.�Ci7���}��������p���ʐ[���p��k؞&;szq�]��V��y������qq��/�D�d��91T�}�����©�9p��C���
��>)���^,NQ�7Jf�ˊ�Ϻ҈���[����~�ڟ����\�l�k�N�<��	��q����㙮��/�\�J�cQ�6�=T�]��[n�&DSL�L��|t��w�֟i@7`�;��`d�ٮ��>.3S�+uk|���>#īO<t��k�/��
����dd��l4DP���hB�`*�w�|����{-��kU��تŗQ�.w��y<�2쁫;�-`7�F �O^?�y�NF{���)��t�3��kAf^H���4��o�-�ђ�U{`�b��$=ѳ�Z���f�iC�Vw�x��g/���a�!̥\���R �����$�A�������
]g-t�8�j�B��G���sEv+�+�|6I�rq+g�����5���S+o��_J{��KQ̑s���{)7a?FAAmv7m�H���Hm?_%��p�XBO�EL�|�H���}%��v�E�Nc��#�8l�B���_�Wu4
nܮ|��rE�מ[���:��������8T�n��_v���T?O�O,7��)��).��(d5���D��g�F7�a��ZD�`�1A�>\�Y���>��̚ �{]9Mg 7N���>� ��0#��t�U���,�D���9�"!�n��?�3�ָ].ඏ��X�z�n����;k�K��SGW��E|���?�"���������J��#h��I�$6�NK�m��^��s�UL{��C2d�F��OYT�t,�}N`�j��t�2�]_��[N%�<�b*��1���u�/�mFi*�#�=,�V����*���`�8�����b:DD�%����b�9�5�qn%�ޗ���=����g2IW��R燖�i���Δ��s|�璲Wx��� 2q��ս�@��{��;�<�7P�:��8D@Q�$�ɲ�G(��h��8VK��m=]�Zi��m$e8�h�5�&��f�oov�p؇���m4�*����n\ZI��OpD��G���0'#]tg��FݶI�P��)���q��u���[<��Bu��Xɉ����pз�*t������ם��4��+�{�k~w�>ڢ8O�7�k0�e���%x+p,P!�~l6Ua�8����<M����y4�^O��P��pA��pX7��+��ɛ7�v�Cf�2����遶^�ѻ��{�'a})�1A��62�����S�ow)�2K��/8�A �_���+�~�9�pN��6��@���4��R�52-�]�&��E�A7�OL1i9�74���%����ø�ҧ!�Z�3��>�V�����	?��=����C��fK�aJ}�4��$��'~�����+s9r��֮h�8i{��c��zl��;�L���,�� �:�ם�1�\�+����//��5Ϊn�T�w�?
9�[�)���!9ٌ����A����p��l�_o�־��������wk���3��|�������"��$d琟'���ڔ��
(T&)b�����2)�HI^r�'�y��|f'��T���M�}�4��E�!J~x�u���.�=�ޝ���`�}C32�X�>�ʓ6ga��şJ��I,百!�sDn�
��Z�K'�����o��,�1��Ý�
�_{��TX�m��s�6�7^��"w���^��!�I�J؂#�KM�(��z����Ǌ5�<2�D��j��=6���><k� VX��귅�l��i"��O"$�R ^F]�1�(Rw��C8���τ��I7Vvd��R+�2"�y�eρaȷF�]rG
�]A#0�j����^D�h�;�O�b�����qbY�`�(F�'�Ũ��I̞=��?�Ԭ0�r�2���جW6uņ�e}�v(&�7�.����(Ů*��䖾��A���\~['3�s��Y_����L^A��)3��R�hA����0�$��`l��q�����Q$�O�ۛ��f٢#�&�E�Aq1)0	M]��gf�J�a���QM������y����������m^��b���P��7�2�t�(H?n\�����-`�yn��وXep�u�[B�1V�s2 �D-����D�fX��2�V6��SS!W鮭�"��RpE̲��l0I��kH̗�ƨ��%�"�8YY���/�����@�n�3�S�mwA���=7A��饺Q�������`b�&�]��^\x��2-��F80�Tl���	��|	N���G3�,�[�]bh�K��?�N�fs �H��ҷ��<1�B5tҵ���v�c=d[ɕ�7p!����&CuB��^�_�UG��ir��Q醴���𤔧K�U{D�D+�ħvҭ2��K�ϋ� l�F<祛�ծKuW!L�m��u �;v���Z����M�:���k�߷��V9� o8���C�����K���dVPc��쌄q[�<��n�,+?��< GG�`>�3yIKй�&`s����Qϧ�!�;���M�͆5��
���oL(��I��� $��Ȣ�I�Uo�:@��;hܹ�2)�P���khF���f
G��2���/2s6��]�LS�k;�!g.#�d:��NIAB��Rd��)�Ja&#C��hُ���T�:�f�&�_#�#�� Lo�IY�;�B[Y�dϜ����S�S��9������}��P�Jy�.�E[��:6xF�BF&�I/*ﰿOt���1�5"
 ���%�Y=g~���B���$j���'��E�ת|S�a�l�v���d&V�����雼��F����ӅW=�΃���~�i���#�zl��)#�F�K��Qhf���O� ��"����<�`:;K���>�INK�p�i��Ͷ�zm�ù������{�m�X��}��k&0�)j[�L�0f�<���ǚ����NG�n��ə�h�y�[�2�
��嬙s����(r��H�z4�s`!�P�M�Q.Ž&�=�[�~}ӎ�kg/�':+�M��sĽ�l
�����ӲaZy&�B�*ET0���4��� �UZ/��Ißn����M��u����^(�1�&~�e��@2睟��\��*�W<���Q}'tL�f&J��</P�7�Do����vq���y�hM�C��8_��j^��f)󶜫S��:ǆ�"`���.Ef�鈖S�h�^hͬ��x�����{��I��W��0��#���٫ڽC�W� ��� ��=��>��m���;�'�+U=� .����g,�����|7����-V�a�=EU3[�=�B`^�[X��G�N�uʧ;")iƥG���(O~7oG�W�r^ss��t��C��|�b�q����E�q>++���:V��j�G��v�51�����s��]�nT��*��B�GSF�GAȬ�Wئ�l��KC���a�[&���x��H�ov�FQh�caC�D��>��&e噦5�&f��m[Q�"��o�F�����>���$4VD��#Õ�wo���S �m�Ċ�����x#�
l���h�`a�0�&ح�T�B�Rا�X��`�s�g�Qȅ���S{��$���u���e�J!_��?*�q/�T���M�b�B��^79�4�0����P�=��PE!�'���Ua^Rk����-��'���v���?��\X��]�~�#���E@�C��ƭ��H�������p$��}�T6��
��q������&>K��`�����0��r�f�����t��@?]��2�o���<�E��}�?��ڊW=��S:k�v<�"&ա�Y�qήi��Fd`�/�ͪ�G�~� ,�f�h��2��+ ��(��<����>�=���Q��_����ޙ$qv�ǋʿV��"�3P?K�ct�� �A�4��JoVW0+��}SC*��׼e����%Ī��ͧ<ͨ��:���$���k<Q��8:u���s�.�1w$�$�� �@��a�nV(���p���,Ζ�w�R�ێ��<�rh����ؽ�5�(g�}*�/�u�G96o�9Y���c鋚L�|��`�.��=2�
��rd��qǉ��FO(��2�����pfX��谪�	�Y�� sC��޿�.��o�]GOqXIu~�g)Y8���+��|Chu�1y��c�N����9m�h�U��gВ�86{��M�ς֓��IX����J��ih�x��zfHmn�����%�$Ͻ���~i���a�� ����Z�f���X�Ӥʤs\85�N��Ṍ�sYE�cu�:��0(�F�
�ge��D���l�6�☬�����!0�|���e,ҤAQ4�\k�m=�q�D�,���&"���;�JS^99,p���p��K�9�� 'j�
�k}Xn�J���g��WA�C��6���nt�Y�A�bNO7���)�3n�>���+R�96��:z�%�}��y�v_M���$b�*,+o^��U��U2��4Yϣ����4P�z��y7D��X*'mus)�d~�_`�(73`=� �n�����(���ں�����'P��t�酟�Ck��@��@~DN���8Y���^8]/���X�4.p����$�)Mc�zb�သ`oT(�m�G���S�I�l|B�2l���M*�D-,����%�
�%��iJ� ~	�����"�<`B�_��ڢa�"�غ���L��+�Q��$������Ǆ���{}�K�� �!Y̾�֪�h��2��{����[����x�6�ҲBO���^d�J��x_pB��Nh��I��	�N�֞����s3�� �^�h�q4�b5�G�w$�B2�ȏF�h�IJ�����{}R�@_=N3����)��z��j�dѸ��(�iUΌ����a(MT��J�'�̂�:7��(A�}ᯁ���P~"��%�J�Ky���mP����xJk*K��lF�E�p�@}�1�5� �|���I�0�?#�'�7^�0hFJ��΅�T]Հ�Ej*��5L�#����*��gAME�jN�0�O<$GБ]�YĬ� � �՚eS�W�^,8!�r�ڮ�r<(�.�/�3��.�?�i�k�1:����n���A`��٢d�C,���bu����n@4��1������O�^�3Puy�x�����1�ӞѾ��ђA[��`VYP������]����?qа�?��ʧ�:=�$�<
^C>%i��<圳=�{rʏM[[�4���U:����z�*�s��e���J�����YN�*�G�U�|�</�U��b�w��QyQ��
F�η'8U�І�Ո�o�0,�e�6��C�cIkD��$���ّb-�`�^��ӶU`��E���K)�E��tE.��^s��h�P��D����y6��l(8��Ԩ��r�S9����~�7��/L�ﴀmH�9`�j�����i����	��"���S�7�\��"^�ZIu�?4I9;S<�J;z�W��U�U�4D�=:����6�UWO�����"X̀��GN��
�x���4/�*������Kb�v}��K�T_OӃ�Cc.R�0������J���`a��:|�c+D���,1�,���WT�����u���r�E%5� 7���YE��T��3�P0�cW���pe��S(�b@+C�mKŻ����J�8����p�ذq>?_�������%�+�6�݌�}�DM��2)���K�%�]Jj�&��R%�gg�[�ѡ�	��D��uhnWP:������B��:�%4D�YN���d�\Xj�����=Ʉ�b�̌�I_�S�ߙ�)��*�Z�PUgPs�f}�̉9GQ�N�м�(l���<�b&'|>���z�E):E8?�?��M���c�N���.U(nv�Ƽ͔w�	�̫��DR����t��]~�H���w�����'��&I�=�)��Y��@�m��c��0"��_Swb>z[������v�|��ËlEWά�\�����0���!��']�|&+g�y}�sA;G*�:���4�/���l���M�0����3J��R<���+�ft=�)1,9��M:!)��4���5=|�MQ9��iB�?%l�ө#s�<!�)�g��fu�����́�R5��~����p-f�"Y�j��]�]q]���PZ-p|�j�*�Mh��{��%�����JlZY����L���_�y���$�<�_a���Xa�>�3�"`��3��ڳ~��$����k��$�����C|�Z�1��Q�~$h����%!�Z7��ac˒������b���r�{Q�՟ܣ���Q�\��^/3x�T�B@mC��a��`#�\fiK�:vz��=z�����ey���r���i���)/�05s|l7.���v�U��2���ʎ�J��=rnǭXv�;���^�P�G�N���N�$��f/�x�87�{�l?\�h����hDڀ�+sh�Su��X��y�i�
2��O��Ƭ���\j��ڎ�30�Y��#t�ī3��V��7b�����=�0�y���~Ti�u�z����[S��ڠ�)���={R)���;��-�F[w��[�RLuV�W��H��T>np�>b��c^:%mSȡy�8qǵ�!�^�]e3�W�Y����EɎ�燾�1��	h� =���D�A�.�i��F->_R�����.^�:�.������VdݨH�h{-��]ɯ���������ƻ?��J���z5OK��y	\H�8�gSO�O;(���1OtGH�:�nn�Jxۈ�)�=w�F��7{���CfT�|��tK���s�Zgk�8��o��jb���!%�AVg�������d��O��g���f��&N���w�
^�$�;~�!�=z{���(� �7��h�{���e���}�<�79e������j�.+;�\�T"4m�|B���/�%ri�h�r�A)Ş�'W��Q���q)IW[�%~P�����iL�U���Q��/�=*���$sE}��t������k4}�W>�}��҈�����
��ʚ|ֲ�,���}� $�<0������i,�,7�b���وO?"<k�RH�6FoO<�4tͫ���4G�9�l���tB�U#��ڥ����_���eG��Ԭl�����a@.�A���.����g��1W?ߵ4�Y�xroďy��P�9�9P��w�msbm�xr5��l�����U�
��4.�:z[�s�})`1�(�32V��'?���!�WmK�%&�g�<63-��m�S5�6��|�ӗ@��Ds�e�G;=���^�o.^���[G�g+O]��jBV�h笈�N��p�F���5�N{>XEٿ���X4h�d@�uՀ���?<Q��g�L��Ҥ�H��5�o=���)|�h�j��m��;O6��|-XC�����j��}�8���
�J�U��a�� � O:w���Ȓe�����x�4�Xn���0��w��Җ�q���P�@�L�7]�����3�����f6����"�M,n�z�k�fY7�t�����4(�����d��|� �Y��Yy���lN%�;�@ �&�M�D0]�*8���!����z+�"�2�ɒ{�.ۗ��	Ԓ%8��#�:�a�{��r�9~Ԩғ�Ic7�`�	���!R��F�J�R�5���Z���A��w��a����C��U��S�����|�M�����f ���W򆍃�暌f�.ݓ��-��x����f���r*��n6£�!���Ս@���*ߡ��F3ܩȯ3��[۴~���Dw���YP�ہu2��'����PM�i1Y���V��"<ϳ�׎��þ��j�3�]�γn��.o�W��$v��e��Q�N�ؗ�t(�g����C����D����Mt���#���k�� Dg~�w[|G&i`���lEj��:���YI��$���pp����6�7����a��aH�4R �N�������𮅰��s�xv�q���	��J"Jp�VM�MBNN	b�u_���Ҽ���wv=#��l�۩�*�@"/o�U|xJ�{t��������di�0�	9y��� {[$璺4 �������p���{@E�.t��Q#V�(TDF�����O�T�҆�],�gY�,j��HQ�KP;�6vcd����Q�ݮ�4M�;�`�=4���nrń�eJ%� ٚ#�Ů�h���I>3x�g/�p[C�ݟ0,T�am����Q�k�K� ���;��"ּoRBl�D
R\!���.�>FrU�����.��C@e�(��/ @XWH?Q�O���u�8�������c)Jq`[�Iڊ�>��ǩ�/���1�����%v�����ez�n"�����PN���C���>�`vV�4W�:̔�g\C��'��T�VwPR�r�>��'���8�V H�ܕ���$= z������4�Y^ׯ	S/"��乁��Oũw!5	K���R:��9IЬ�$Yu�<�c��:�0"1����w�*\���{n�u�y?R? �emYP<A,�p���ۏk��]�P"���gW~��1���r���*C�I�ҌF/�,㽝i�Y��̎�W(��,����ِ(�֚E�������$�)S��M̯b_�ib�U���x%kj"v�F����x͉<�����b���w1��〪eb^���k�-%��M.�+�!��E�����KҴF���x�R���y��;����Vpx��E��l�|lC{@���n�G�S�{r��t��b�W�,F��J��Nb�!+UU��
�vM�TY��41�&��1W�6��I4#��l��e�.O���dc6�����t���^��V�I�-�=K�7B<�i��@&H�:�0}��|�w+������z*�m�䯄��`����7L���E�-Qk6�3���Z_ƚ��	�y��[����� X�@=3宆`�e�ä� n��u��`c��"S�ȱ�<E��x{��0j]����E�w��[�m=U���MY	Q���|h$ ���<��Z�G0@�׀�7��\�ӊ ��,���4w��N�<���[�W!b��/Q(т٣�t\}$R�N���Eѿ�4�W`��E��L?u�,���&@*	�#	��i"I�_�D�$��/�';#V��U��q�=�M���4��ӎT������@Ƭ<�7P[��2
��r���θ��sL�ӂ��f�AC�,~iI¢�_W��W}G^`RE�K4y3!F����.�%��)�n�I3�!M1u�Yj�l�q���s����i��>����y�mؙ�?w���P�Xxx�c]�흸���X3EHB��^��2A�
,�\U�A���.��fI�����D�b�zW�cP����×���<@�ܙr���Qt��Wft��`y�&
����Ę��0E_A
 ,f�r��B���~4u{��i.���d!F�r���K���?{�	۠�USV��q�g�c�f[�1�
�j���E�L�dZ�W��9�?pQ������u����U�j���܄<oL�#w7�I�?3s諑��p��g��BL��9e{!UO[n� A1�{��j��-!3(23d��
�EX���3���&u~�cC����eSz�o� d�`��Anz[yz�'%�"1��^�QHxyQ��eȐ�R�6�҇ ҽb�,2]J�g�^0�������r�ֲq::\�Cx�� U�{J���
�Q���.uY�
*Z���a<�*��u�r�U�N����T�p��,|#JS,��mzin��H�'�� U`V��&D��t��=����#��н��nK;�:x8�i�г5-GbZy*
��م�Me}�K^����萳�aS�(/x�31ٿ�]$����D7�X�`u���|���u�)��y�rkO��{�2o�aRB�����de�����e��$*��/3,qB��9�'�� W��?
�B#:�d��Q\('-�e&^m1�M���\�CJ�4�K�d �=<�f6�M��9G-p4�W6�8延bm��u���А=~�O�M����rt��b�4+=�<��GP�E]��J���k�WG�7�P�*��XM�Ⱦ����A�n��Mw�ְR
��,�1�����}�����&z����Y����X��{(��O�xL������&�4R�@a5L�2��k���ã��h�q]� �����}ۨ�"��~�����m�٘��B�@��!�xgڌca�I=�üvP��o-�zp�?�ByA��&p�� _^d=ousZ���(tS�<r�Z�5�Zp���jc�������>8y��iڜx+m/�u~��m�/�F�0��P/͎�M�.����y�q����v�_+����Vs�܊i�&K��2�(:/zno���ؤ}q�\�-���v%�k��7'�H�^�q�0&7M&�h�pe�A5�	��Um�_n���<�>|&/R�x>���L�a�u�!�EZl��﹃mnV�,QNQ�}ӝ�����.D5/O�/FD5Ά��e.�H6��A=�If݅`i���<�ϱ
�J��p���p<dEW�
$���[Q�*��l��Rp2$�}2g($.R��j�_�����s�.���+��{	�z��P%����T�t�"D��dorG<��_�K"#���<�.�q�\�|B�cHp\H����%=]���`�q���������������M�?�!���+F�������$k\�oY�x��g�\+Fe	�'l'x�{?�T�ia��i�?~�͒4��~��ˆ z�]t���;���:�U6ڟ�(Z#��c'��(�Őc��I��%�x}R|�k�1��qB�P\��8
@����u�^W'���@CIE� �*�`.�x�$8_y:gaRAvn��,�Z��5F��yk���- ���,�ZF�.V+�,��T��c�'�ֵ3�	�8{�S��رl�v�9��V��X�Ck�5�P�(S�~F'E
+����d?�,v��kTOMXHm�!��.92��F��H�&��"7(d�^my��o\^J�"�%�������MO�f�r�$ʣ2deG�ƈ5LG�{,�Rs�� �\��e� �&/�>v��`ΟQ1Z� `0��}��l����>'f�3��n�7Fv������^G�{�ϝE���x�?�u��~���(c�N�@�j�=�I����Yk�C�X�N�t��m�p��al�nAφk���gd?��r��TK����ݗ�C�����t8\	Q��k;|��u�m%�*��" !=���n�K�,�����$Wӂ���`��g�O<5C?�(N�m hh��Ӈ.��oTH0�oA&�kd�|�ȮGs$�q;N�|5C��%S=x5�}�T%����S�p}����&���A_7OQw�#�.W�2��E�װ]2h�	S��=�95z���-�E�X�m���Gюo�}�ZR�<C��
:{#��]�����@7ij�伅o���	㰢l'MP2��Q>�6x6�n��vs+JL�ء�0;}��J���rz��Fa�v���t����Ǌ��,'�(��09�n
��f�������ߧl�Z�T?A�f�<�W��n�pl�x#�+ȴ"	�0`��0�#���e���gWq]��	v@ꮹ��+h����5��"��-��I���t��qr�;����cb+��.�G���Y�ލ�M�$��x( ���l�1����rF�@I#>�<pA�	E�6�Ƴ��k�L���u��*�E �ю�����a^A�s�ؐ����2��"���EP,Z�e������ъ/5v�`�5�;zz��W�	+�v����a�M�/3چ�+ۜ7���)��T��FVEkG���P��۾�e}t���3Ӧllҟ�;�?��C�l��o��3[��
dl$B���1�?;۶N�.<��t���7��2�A�ȕA��zb c��m	�Ы�h�	���V��t�a/�,�x��d̒S@a�@~OǺ�*����L7��?�BZB�����%�ۧ|�}���S/�J�/3Lp�'|��0����������j��%QM��4�ۛ�'�7O���@�E�3���J����g�*+�m�0q�㶙t?��>�x���)�K��]y�Z��C��^a�X��23ݑO�����A�Q�x<���S��@a����ŝPԁ�&a/�$sy�7؁�h�t|6"	D-�r�oH�r�����ī��-�[�i�N� {ko{@��n�'��J��U�?�Pk�@j���L�����F� ���)3!QO���o1��d��'V�Ӱ>L���X�B!�I�O��b�Rk����2��#��o#��P�KCd:Nm<n�Q#���D;��.��)z��S滼ܺ)|l"ĩO��*����=�a�?��k�@F���m���2��\轁��sf���L������_R{$J���v��(�Y@���ʤN��}���mL�k�CǍͻ��5<�]hj{.D�ֺh�7ٰ)Z��}U�'�>S����z��q$��T���$m�Ǫ9d�h��+0��� e��9�'����P��1:S<�	J؄��l0����T��1Hi�Ǳ�� �9���A���@����0bz5iy��QN�'�ѻl�q�L�΍�A'ri�li���"{���[oܕ_̧�v�T,��Ƌ���3�y(6�:R��ER�IWrl�����oe�^�8�Y%*WJ;a�ɝc!J��It_�.x:����F�W-�,�=�Ut���L|u��?�o�X��P@�D��jXEq�S�	"똠�K���K�z	PP�s�}g�_�+%��1Y��SG��Ƽ�b�!��Z���R�O,���V9��!�m�����x��=I�dWRHz�n�V�#1���n�k���).#%���Q�`Cw!���oϮT^6��8,�|�t�%=8���[V�w��<9*� �<9��)i����W�'Ɂ�'-�}[o�F�!��'��p�j���:�J�`�\�O4sbr�4N�kO�t�xc�y*�]^5��`M�J6�a��X��́bQc1���#�!��� �����F�Iv|L�"͙����M��K�w��&��bU�4�R�"~�-
�Be�i��b���י��{����R޼�G`�iN�U�ն�>@2��L��[� ����,�o�-=M(9P� ��o����HŲ�\� ��M�x��9���*�h��_OtQ�M���ڀ�aF8�����TQ@��0��;���R,�12�2����VB���%pX��4'�FuɼI���0
X�����`+���PS6�&��*�~|!�S�.b��g4 ��&7+;pĔSB5莀b;�K!� s;0�y	�3������2V%�B��3�O�Kţ�t���N��\55$�ޝܵ"�Ǖ�5����Aw���mwK��cl����o��H����/� ��H�W�
����@�m����E���?!��]��2��t�S��5"�S�M��ܗg�x2[�ǀ_�����~?p70H$Kl���������H_��I��� WD���P�á��	�l�g�u�1N'r�&"�~2�X@N�!
�ԯ�N�s_�i��B�.lÖ�1���ڛ	_RkE����0��W
��O�������,�Ӗ�K2�1DM$��*n`զ����
����톟���g�������7�-g8ћ
��Z��"��t���n�� *������֗��[&��B�����@@Ep�}��e��x�tԟk�f��!��J�Nz������X�_E�"Jّ����J�5 9Y��L��ǻ�w��[�m���3sh���M0���%�1�o1�{b	U����G�퇫#��밝��5X;�U�@���Kp>�w?�["w��Wu��w
֍�������q4�V�<^������?�N`	L�G�v�ٍ���x=H��5=�L���㟦���͒�y�����M�&�H��F��vt��%#X�P����]>/MJN��!�fh�Y��(��T���L.�B����ל������ÀiVf�m%��'��IJ�~!Þ�:čk],�k��_�*�T6"��x�0O-/ܷ��ﳪ�۫��^� V|��u�|WL�aLl�����\Э�)7i ��.#X�q�K�*!Jn��_4x$����a�KӼ����� �EZ_������3�;���-"]%��$>�{�S���������߳�/�s�l1���JL�����3[��;�>�Q��������z�j�����������#_S�{��o��T/ΰp*9���q-W)��D4�(]v3�-��~Ϧ�6Pkq{'f� *RS�E4&j����-�vZ�{��hf��N+(_F�:��?Qo��*�m��)+��΂��i�:,7�oj�ڔ	Ԍ&ٸ��7b�4 �����ϡT!3a�w��:��,���ȴ����k;�U�bFuZ�NYP����+��O�Ӭ��!�m�^���MCTuy���B8 ���\��+xfk�Wj��]T�O
���T�0��L B��
�I�Z_)X2"�����[D�$������?�u�Wî\�@`E{K�6 :h�R]�D�~����$e;ފ�rB= ��;_�{_Pk��g��d��d��61�aK��f�.��<Rr�kk�|[���/�	(��TF'3��Q���룲�i�"/��`����Dv߇2z��?,w@�������n-�M(��Am�q`��_iV�����(��r)#,�D��9!�m>�[�Z�_��]AM
��3lq�n2�F��u�I�@5�iV9B�AX�A1�PRd!�Y?D��F>~3�6�M�`,�i��`6��!<\F3E�����[�K�\ f����$#�0�HT��Jo�4wWd��c㝟�Ϸ�q^8%���+b�3����� �*��Mz���ʋ�E]G`<���
�^Kti��-!���#�:�6��yg����|usi�,>�������`us��Q,�HtA�~Q�4h��S�)���
�9R���z��(�/Ֆ�ڇԤ́ԣ��*T@@����7<�
<�v��<N7_9{��
f�m1�b�7��o¢��*RI�-?�����q�� �[R���'M�$��z�S��O�ppi�������yk@G��bjÒ�ƍ�1M��[����O5wn��}���g��ѫ��3qI��k�s"'e��&��;�#h�����$�2�-˼s���
��wanO�e�b޳ '=�����9 4����j>T>�ɯ,!�34�[A�����M�,��&?�ɓl-��������*-���y=�U˔�>��M�d([I�����x�C�*�"A=^���w+?7�Zf�O}�ZS��P��Ytg�P�dk� �Y/�	3��A�����ce*�>�������3�2e�o ������6��_�k�����/���kD�8{�'é2^���ϑ�"BX�͚��������C; �#�����$gD�b��+��G��A�1a��>zyTMP/a\�2뱜�ǳ�:坔�����	1ç�����e�9]e��6V�x�Zv�K��h�|Y/~��@>Y,Z����fň���\�]�#kX�
�!���*�3\3Fl��w��<�^�E%������6iV��^"il��G�8�D�@�ӏq���e4r�o���Rl� ���~���Up���KT��D�M*�<w}<�(DѺ��V�uC��5�*0��韎�VzE���L���x���\�<��^�oo��z3��t��*E��,d�0�a�F�aV��*�'��Q���Q�ftޒ����F�ѳ��1BpY6�I��qy�|�t�~��`<fNSZ�z�����ۂP�\�U�=���m���7+��9tE��:],�w��a>�2b�pDL��rO��+�	���wW_Wd�+X�*�T�mr�c*b�}�����d�b��S��ta�(a�E�֍��)�r+`�S�`k�^��;/���ը=.�:��A�k�_�O	�����8�X�K���s��	9������?!�2g/CW��(�3��L��!���F��r3�"ѣia$N�ˉ��p	�I�-�`�=Y3��R��w�4�����;Q�e��oܽr��޽��CI*Ι�TN���X�YhR�<������;3e��r����T����������Wa2�vxonں*/��ѐ����A��
���a(� ��E�&����(���+Ԇm�� w?E@��
?�)MZ�ht�P}a�`�6τڬ�W)�4��@�)���5�ȸ�������D�:0��r��j	U������8�i�MZR��?|�]��&`� ΂���a0;��A�G��	��Y~���$��3pИ����=	lK�V0�}�`g����h�1��Ë#��v��G���j�i��nz��ϲ���� �K���!�,�K$�qt��p�����V�_�>&�϶G�̓U�]v<�y��篵�ƒ�������&�=L�O�$�c�麲Xz�JX���`�賈j3;�1��\�v>Q�Ւ��1ό�?)��p��Q�.ʁ;^���a����� ��g0����������T��H�A�"|�W��<�b2�hO<[����%�$��N�6�����D���E$�C�-�xDA3��(��Ϊ�b~�S�ݷ���7��� ��@���s�q\��h��3+�R�srgST�0�:�U^��������Z�����N�#�n�0G���B)y� �����/�$�WA�_o��@=�-��C��jG�9��r�\$�(��$#d���H���R�K��i_�E ���,�Ix��d�:/�F�eSsЙ`4��I�?��`��F������g�S��y��r�������]��w<�θF�����KN(�*�"gݨm|w�!�S�4��d��呈b,� �t�e���$B��|�ɀ!4�|�>�p�����v�l�o��k����eݮ�wW��d� $�s���0��II
3_�g������veq�d{�4<�3){�=n�{��\ʨ��:�	a0};ۃ8ܻ�'O2i���hu%��S���6F�9-����v��$���B��gs���Ί0�I��n����̺�`�_��6��R_d����:9 1#����x�0w��H6/1�qʆ�]a�};߭����a����j��Ԛp�i+�B���2�Qi�60M�'f�����1�
�^��m�2A^���p���Z�D�@�D�p��K��
�{]E�������X��W(�3ڜa4����EB�i���ؼ:��Ҽ��t�Q~l���p�m<n�`L@�%WF��u���������܅S�(x���{�
����5���x��&b}j?�#��ƙ98������I-Ɩ�*��A=��v�X?���[�FP�nG��F�_�.;G�z�'Rcp�40wY�����-�1�-���u�TU�I���W7K��,�9�'Ze6�Tq� ��jK�Q-Q��}�"�5�kd�m^D���!�؛y��_<鄵��n����Ǻ8�m��|�� U�����[���us���0��ƾ��s� �Z�����g����ޗ��Դy _��;�h��C�\f��O�4��\{c�r㬁�1 G���Ύ��?+���0é~u^@�R�;�@@���a%T���a�����M�\>����O��-�F*H�~���}���-RRP`�z��7��n��8�w!<zC��xB�L�: @���B���f�Q��!|�n�r����c>ݬ����U��-k�ϧ���L�^���ēG�����'ڜq< ��GbQ�<K6ic[��3�Z�I�N�D���M(�X��/i3}�����os��7��z���nR):M�6�?v� �9p�AS"���zev����o4=���= ����M�w��I*5���K�Ox��[��|��C��F3�F�0�̹�-q�cke���M[oV;h�sސ��x�xx*����I���yeUn�.�8)�{�.A���|:��M�w/����d�d F7ޝϒ�\�|���2p�Ym� �^:�wG��$�T@��i͖��c��S𙂙���O�S+vt��u�<�2�-�n����1���[��=M�p����ѕ6=²9�y2m�<�������l�B1���3"!i��=i�y}Ӫ,�/U��d`��5߇�R��,R�7!=��P��a�E.D�Gn�� �%fJ�D)��G��/)@�֞� �z��-��kb����	xbF>U}�<5)b�����/5��^�X�Ɋ���]��	�ϮG��*���h��~$��x<�U��N�2Y�����KA��q:�4{�#�=.R��sl��S<		�E�U��^hx����i�'_�֖G늶��ͮ��Ȱb~��d�N�\#��b��P__Ќz���K�]3���3 �M�ד�݋=m���OO��݅\="����_��͸&�F�n-��
��Ҥ0�`���ꖛl�r%ӂ	�{��(��W��%Lx��>�q���k�z ܳ�F�;�S4�:4�!�QS�)��R#;��[Jk&��Ds�6WP�ejeU��\ə��Cp�_!��gU��p��+*��w%ܜ�Jܦ�f&�rC=���+׽p҂����]K�)�i,*Pi�\�L���	�$s�ۖ�5_S�n��)�'b����k�o"�Ye�[Bl����1�Z�T�_�)�` �9���4�{�j���\O>8%LO�c�~�J{N>�F1E���j�ETZ`�C�K��aK�,���/�J}sCj�D���
��N\i��F���>�m�_]�է�����7B*On�6YVj��9����Q�q���/��GDF��E��f絔s�����Bq�͘�)��0��ֵ��I��&S9ڿ���(�<D9��t�7´�9���|:�_��gr8���%��_��i먠�ؙ�%1$�@`�����?�(=q^}�0VO������red����b9�gkO��u�	��ѕ�LF�S���!A�t��4�#D rBE�|S�@dG�V���1�%�]W^�og�I/@��Z����e�?����+�n����d�D�k7|��p��b:7��8%�J��»x���\�-��&��*�ҽc;�G�_q�2��&�_�q\�ks$�MuE�Z�7���Ŏ_�b�bs�
�\����bW��h5}!����=��;r5bk�Z�S�z���C�?[tF:����;���8��o^1B�����&U����Ҕ")(���[v�r���K���5Ε"2��%c}Z��*N�A��5h"u���u���|{�n�����A���gDe�̠��w�Zk�[��^����a�.��OWw���ė_p�yG?�� kf^����vxܳ�Rn��d"\̂SJ?�ש��l����#��J��8�%��+c�h3����jh��-��q�f���'�VL�LU5�BFA4LC�3\�b��1��!+�o�Sc����{а��"�_8�c���ʏ�T��C*@ăk��CD�:}f�g9��� �jbB�MT���#���r6澗�A_�r�j
�{���s���i0�@J�:������ ����bP8!^���G�=E���Z�U�U�G#!��a��D/�>��(/W��(9	Dy�+}���N�z|/Y+����Yd�$���g�2U�w~M˛f��}�^tf51�H��Sve���%"SR)y�UB��e���j��ї��2I_BK3/:mã�> ��"�[��"�R���-��>����;B�+nƠq�KjC1���\cߐ����r�Z��i}3�D�6^Kh�,�ǆoi�<l����T]x6OY�'+XE����LP*��3��=� ����j򉄚�]n�ֹ��$��k�!��ת͊�z���x�Y�TӘ�ṕ����P�� F��j[<3�X�O�Z`�'�$?�}�4��W�P���W�IFx�.g�����$��0�Bm�1ڱ�᧳(Fx�)j
>�;��[h\�`���	��a��(���!]3�@�����]�ԩ�v=����!Q��"��ql�?�V�)}��Ɨ@�WU��}�Sz�dkn��Jf�԰<8I�H�w�)�v��Aj��BON�~H��k�U�(�P��8$�K[��t=�y� �x$����d�M�#�PFɌ����h�O���2����C�2��B?=
U��=~�0�mAS P�q^$Vڨvg�H|��tǗ{�<����0f9"傼�G�u��h�R���xH#`�Ή]SI���?ep{�B�@*串����:*�\�҃��S����6p�v�!y�t���^�����(,��$��E��h_��F�����栊���eg"�^Uj�h\d"�r~}2�i3�Yq�3'qև=���N��R0Z�X�^ JLˊ���Ƹ�K������%��}b,�'�&��E��<����݋{�
}n  ��D�cn��S�vC��02�cc���p��X��K��_�r�J%���$��CK�N��ѣ��6	��]��D�߲��Þ�S���C�R�:���J`Zmc���AE�����qx��T�ФM�,㯪�����5����.���t�-\�roưֿ��X����uWP�<�O6�ٮdNt%�
����F	�&���̒(�7��W�ތ,\zM+St���;��"���]s����)�7W��[4��S�~�t��e��^"��
�(q��Q=f�4d�9�@�O�]l�����o�Rø�z�OM^qI68�����,�_����钢ikÚyHF2#^��~C"��t�/N�Wц�=�\�,(Q�v�>d"j�d���d��7��>j�Q�&\�1;r���+��n^��cT�
���@�����Q�1(~8Wf	eIrp�������&O��M�&(�Q�kmߵ|����<��~�a�'�� ������Fq��J\1�Hǻ�h�=w�"z���[2_����,.~�\֜g�&�?���j��*�,i8bR�B{l�ߞ�X�~�0�v�gr�2�Q]�yn\jvJ�v�h�f���]��2~��d&Ad0g+�?/�;��2Lzq�L��`Ѻ�]�@ "�њpBXr\�{n�˅s>��Lԏ�G���:l=Z2�р�G6�>�Ĕ�k��Ԋ�*���l�����)�z��K0��SA�J�����D�X�V�9Edb*���HԖLZ~�e�S��X'��M�ee�w	�ՏԢ���^&ww��cs}�mX��m͈G����8��G���kXfMRxߖ���|8�Qh]�,���$��O��Rl��p)��=PL� �P���JD��A�W���nڙ_GNҴ�d�ʦiS����(ڣ�"݋�&��FAVR��'
���pD��!ޮ�.����k8�"�/�Щ�����Uz��"����2��n@����Y����Hع0^�A�{g�X��`e�.C|�	�,P?�~$M���%멢4����B2O=Y���DPjm��w?_��-)��멡.�>o"��i�>�*5%V/#tBil�t�zډ�f�j�S�v	�*1�A2���8i6
 _���8.�Sb<8������;�JC��j�i�)����m�ȧ@�Y�,���,R0���u�t�'�F\���>S]�1c*�NIl�������>����luC�*#A*���A�Z���i�G_@N��~ecdQ̅Ae܇�8z$�[2gl���H��!M�q��^C�Jɱ0���'���0��Fyd������SǮHKT���ae0�)�,�׫>#�~����>QR~�x�;�+�W�|�։�v�\�<L�����:�+�@,rb3Y���� �R�I������2���a�ί���K�o+�����Ǫ�� -���BF�r�9��� ��}��̥�\�I�W��9��XP��T���A�<.�����*��^����նI�Qb�����	�1n!��f����@���DR���"�_�n��߿�^~u���إ���9�إ7��gƙvh�n ����~�ߩ�M?l�車�s�B��9�~rXc�eI����VKH(_��Ym�dH�:���KKq���"�����ZP̘$�/-k��}x=Yrs����2F�����<���y��E��<K���i�Z��X�J�'�}��+|/V:��Usђ�IVP���O�B�?��{@%��E�n��_�[W� �f�qaO%Gߘ�Q*RL�t����W��1�0ꕫ����6�>՟��-����A�(!��wr8��!����U�䍽�<j53�%ٖ���;^��j�+ �2g:���!<}<�i1��cU��wv�����!�,��2{�q'/�$>7>j�zL4,X6�Vzڡָ7� N^~E��(%���˴�����R�=
]�^Hbq'�!���3f�s��0h��%��{�?1�M$�#��G��cC���f۝q�/,@(��]oTe�y�/w��&�<_���w�wl7�q�,j_�m8+B�'���Ț7��%�\�Ҹ�|�!3�{}�d�I�$:$�Yy���I1 MK���</���l�������KYh2U��kE)�1
J�sμ耤J@|[����ZL�R�oBS5'σ{nI�d�rtՋ�������ZV��G6��8'���p�'�j/X8�l"�&��{�c<��ep��_U�(!K^�����.	��\f��)�'Dp�����+i��[����J�� G�UB�<�hLoU�t�S�e�Cȸ}�'�7�ug��%���_��v9.l������<����f�3�����X5i ��,�4b�b��$������+���:d2o�/s��������fK��{��J\>H�8����������6�E�޺�xM�c��0.�����~3�l�AE'�)y��A�Rsiܯ��E�uj�]�ry�i�¹C���,&]E �q4bϗ�y�]F��"��<��,����l{�"���#�)�t��I�v�0�)���i��y���� ��A|P����ߓ��|o��ȑL9��T�\P]^��U��^k�z�ޗ�K�Y��Q�V�r#N��c0ARi��Z���?.���>�,e�\��Ra��0����yF-)v"�F�7���Jb֣5#�M`�i�書н�P��-����v��.��;4͇l/�mCD��)m����,�v$qE�?������Svmn��&qz@�Z\����޺�w��'?䠠~���E�n5;'pX�;%4@Y����(�V?;�C�d{L����M�zD��K9��~Y���! �v<*�݇���V���o�0~l8��hQ��4Ϭ�sW�@Ug�/��{e�q�Fd<X���o����wG��3��R=�V�]7ͳ�0���G�-(B�n�	������&�ɦK//���:$��NJ�(��)g���� ���x�C�=~�̉���p���<
l����n��D�p�)Y���a�.��$�y���xz��?6������Q�lO�.
�H6�,�����Ǖ.�&����	/���;�Y�)���������ư�5��u8���2(pp��z����4;:�/�9zp��C��;v��
3�9��͕�U(������KAѝfI�<����13��C��^\s� ������&���U��M�����������o��_`��.��H�@�ƈl��]�m�ߙ�r(wi,��R��բY�S�E���˼<O�p%�9���E�=0�X�1qs�=v��d��Ed���oo�����	�g��rNA= 2�CIG��}�_�v�=�<:z�LY���ݻ��#K9�Y���Y���m?`�C�>�2�?p�K�)�	�\q����"�����lW:H �T~o\�~�ǚ�!F��9$�;����uJ���zI<Ë�)����S������H#U9��!� KV��v<���zx�g�q�<^ Y� 1S�V�/3���X�[᭛�W*���+�yJ*�: ���U��eR��=�so���!�M���</�v��D#����-�0[���;$��b��rV��������,7-�W��۫G�b����sC�B�)��i�����<�~=��ʗ�7�t滅}���h�V��/��{ ��a�M!���	�][;�{��}5wgR�I�������'����1=�`�P8Ǻ�UF�@�h��ݰxb>5+Y��?v�,shE�s�R�κ�tS[�A�����Ce]�lu�?��`���b4x��F�8�"�j�E2���ǌM8�� �r��hs�<&�0x�}_���'`ڂ�׫'����
��9w&���d�6b���y�矽��H!�uƑH �����L�_���t�����SX���A��c��Z��#cN���	u4Lۣ�S�{i��g�z�a~L�i��F��D˜Vu�7ժ�%W1�p���M�Y5+���!~$i�4�|�M�t3�3+C�/��^�{��b�i�+_�s^	L- !$���9�ǩיX�w�˃l�wԆ�;G4����u����l�ʡs��{��J��!\wîM�;y�l����a>ȫ�Lhܚ���7�>A�ǀ�R�"�y9D��,;��@���;�*�t�2z�a�1�oP+�:/���6\��C;�PC1<ɉ��WŦ;�%sJ}�s
��%��FuS�M%3,uJ5o�$��tܨt2�sO�ec��ɝ�2u6U/2fb�����kbޑn�)��p�W��'���RK�|����s���N*��0$��V���R��%�ز�	W�{��)V�\k�����v��/\��_��"�s3��?�כA��D/M�@,��5�g)��!��`cٻ�����&r�r^1�Jf�ɧ	�O"^����*�^���	��^AA��L7$@E���Yp'��D���d?�3�0-8;����ʌ_?��?�t�we<n��w��N-Ȍ�)�Y�I�+	�_�̖1qBb{-���*�?���xV4*����N_��)�'(W�R���U&����j��I. ���02_��A-� �����l��&0���bX)�|��DǍl��B+���J(k'j��c�=�;,�G���.d~�~�kva�s�b9Y*mt8�~F�=�CH�`�Vh-�$������m�Z��$LI�++9����ۢ��x�?���w*h��+���Y�5/���дv@���8ŏ�d����-/����Xod����b�!�cM���U���kx[Y��Qr�w�� PC~������J�^��JnU��7,6h�;�ܴ���l���'�!|5�z����fEy�@=%��X)����X�D�3��:7�cNȆ�+y���y�YQ�N!~dV*�z��G�#�S��[w�*��p4��lع�(ܫ(�3�{��v!���I|�s�\�bp6C~�)�j��|��N6T'zA�O��A�#�BQ2�<��\�rk W/���H(�ड़L�Q�ɠ�v�0��G��ߝ�s�gP+�Q�8�n
Sj|�ُpx))~!`�q.`�Sfţ�;�/{�@�o��X�R�={��j�&D����_�+J������o[�/_�hB8���������*��ۥ��K�#�Z$�.�'�IX��_��OS-G�����?���*á']/R���0}x�;cuw���4Pn�ci缉��� �I����+}�P�Y����^�{�ن0tڍ���4V�Н^/R�)��"0$O�G��E�n
�x?vl���s	���b�%���>`*��t��G#�(ct()2���d��O�ɉ+ĂU�Cl��gu�;�5�>H[�
��~I��I� �,��Q�Sus�t,'���Dn�-wKw8�s�R������պ���I��R�I� ���'��BRs[*�� �~Q��{e��TR[�uu�"�1�]c��lF|���F[:�O7���5�)@da�:<.��d�+��vv���y�tXXKw�ݪ<��'p��r��cY�Zx6��FveƘ.��<�:-����.8�E	�����+ݼ��oz����k>�3���p.h{m��8�s�xnד�isdZ��"�J��#�cЀ�ȶ��2\_�	���ʑ������`�WJx��H]�֡��H(A2�e���KwGM�*�3 ս[��b��W�B�ƒ��_�a$���-�P��Ћ�����NP��?���T�����aA�x��!=�d �N�wJR�)L��ɂ<C� �Ŭ����j3 �}2�Jh8G��Y���~�� �-�i��}��
��N�7D�򝞣����cL���r}.�:%�_��ܨ���`�?�������5 �Q���m����/R�I�cƦ�4��`z/��7Bym}<�	�2;�m�6��2D;j`�JZ���Cw�!�9�	�^�IO�p1��.YA�3��߯�%�Ď���\�{����1�W��.O���@6�أ�Ve�z�i\d���9�!9��}M؄��Xy`Rmy���o��0R�l���\�ZG#$/�B+��+R~���t�*�ךa���B���8��g֤�d�����~��P��}&���y�U�a��/�����\� �����"m̩]����S��߰�:{5�:6�2꿙�I� �X�	��D(�8���nq��˔Fԉa2SG��*�n�T�\�m�\��%�� �ľ"��+�ӄ�]ai��	������5�%+��Z�2t䳑C��ߞM��a�K/�ͪ��8�r^vNr���.��Y_���5le�!	�����k�� P���eC��/��Q_�~ݒ�_�>�72G�.�c��ML�'3�{8�: @6��3���G�p��Id�$e}&�|UaZ���`��%��ϺM��!ؓ��Te+�xl&�+M���J+h{��4.���V�4���ԯ�#y@]��+�u�����G��4NF��|����ۑ(��r�i�YF��P��(�߷w8:�(���A!L)�U�4_�T�H� i��s�s!#�OS��̯��˷��h#�����Y@�:��L��kʲ�Y��"���d\���a��������bT�ڤ!7�j��*�)o�o����zഺ2�<�Nk���F������b�hɑmiǱ�H/���q��I�� �����̪���A�$KE����f��"'ቄ��_pB��!�GrO��9�jm� L��Z����xPL��(�]Ӛ�݇Ga�fM��i>�(3��F��6<��ba�,�SDp`�uE�t���Y��*�ԧ%��p�_��?kY_��7�	���Qx�:|�?(	�O��a	��܍��}A� ��DI5"g}k�,iqT1M!{�%��n�R������)M�E�lv��RZ����11�+Ľz5��JX?¶�>VŏA�I���=��˃���]�ou��E���Vj����{a`MT���''*vd�6$R��)�Dh+�p�r$��r$bn8���8�<WS��q'�΢c��7��q�J��h0�(�����&�1!P��ep�S
�\�f��{�5�ZFNU<��@�:>���*���1bn�5�~/,�p!��� �<w�#̭@��J5佈�-<�g�1{?މ�Z�+�b`&`Z�7�
������v��fe�<����w��H��n��RXc�g�����ztEb/�Z��z,��xt*1�U���Ɋ[,f}d,��9J���IW2e��~̝ �2��f��t�&+�LhP�:�C�TNm������ɓ�"Ǣ�P�5L4}�J�@�:}r>>���Ђ��~��C#���$o��*uc�R�oE�L�" �*��[rr��E����o�A�T;����O�E}����z�E�m��JMZq;G3k%m���9��Ix2�\�'���(��2�?~���d�cBzܵ/o��_
A��T!E�/��Sr�"�JL��*륃*�BPÅ���a�$���}1|�Y9�س�;qN��C�l�!uu�<��r��[��s�W�\	���������
�,Ux��+�8�X�3a���jx������a�� �Q>#e��t;m���!~D���5�7��NI'��`�h:cmT�vO8��xWb!�����|oǴ7?-_A,9�kK�W�N��8J��>�׫�j�6Z�^�����)�66�B���x���D)ŗ�f$��fOh�L�Y�)���F@�D���Ǧ��M���Ǚ �R�F)�1x�њRv�%X� �r��w�
A@��e������W-��g
�䩪}��(�,>�`�?`��gB���Hܚ�lxlȺ���p=4�d]�_�G;N����9���9<)�:�kf�k]��#�������Gݞ��	�2X�ì)*}�kڑ��8�m�7?be7����7��̅�����Q���J��@tW������5�;gh���&ʖ`YD�lY�^|	\�'�jS�m3"����']B�[ĸb�����r��S��U�΁KAѻ����`#G��}j��GF�\���ĸLLJN��!�E���N`L��v���2��h��.7�s��[��f�}�ꝶ��_\ ��^%,`��ɾ����ɷ� ���P����c#����	�pe5�q��w��qo���L��E��fFZ�ܳ��:Ϻ��W��P�}����PO�E �{NH֏��a��v`�\���_4"��
���;r���q��o,��t}b�/B��a�WWr�C7�k����~����ʬ~��3\؎����yU+�qm�j��G�A�ÛxR�L�cv��]%��+�*���M��`���:�xp5h���n�����"~k��,.V����1��`cw��Cj�8���2���w{w�g��z3#�����e���Op9�P�I�$.Ĥ3&�M����G�<���4�c҄xfhN�T�^3�L�93�,ѷH�5ԅ��߉='�H{Z��$�!��i)�B��o{#(U�ߗ+w"�X�
m� �v>-�wH��ҵ��}�����k���k6n�V�<���c�(�*�"�%'w7���W���羑�`����`œ��X(j����E�ޅ%����c`� ��$풣��w�o���ݿQGl�n����	�:-�>N/n��=L����qdT5���
4�Z돽N��O��AN�;�|�0��й-A��iOp4k1�~�C������,~�2�GU�(_�╈+����i��S�m=�Z>q�k/@����R���"�0�S��WL��	���'`���^݋�cb_�UeҰ;
]�\�"��T˲�%⣸�P�0�D&A��:��}�c~�8
sJ$�1o�W.��d:?�:虥�2:�h0 ��G6�<�jP��P��,)��:�WN�HG9�AY���Տ���r^�h�b�=�=�
�o�Z����YrЋ�(�`La)9�l��yJ��[�,�ެ�r=�(��a�te�������޾����7�k�N"�h�<�?��eb��{��w���E%6�N)�y4�]5:�Z�&�Ͽ=��6��V���<�d���'������\Е������cޠŉbo�^�Fp�7��P;��g�S��k���oq5�S*�BM����&mA����N_Z�y�uYPM[Fb���u��K>f?��h��3_�\��78�ٔ��+=��e��4:�t�L��x��ĆR�M��9-]����e9��#��Q0<�*�B���*��ֆ�.�[ߍ�b�֢݁-W.}��'�G�T��z�d�*J����j����G��%.�t�X�����p��U�ڪ�H����o���k���+ٖ@2���{;����&<(F��f��v��0,"�U !@JFn;�s�&�@m�EM���ױ9�KIi(�ɒ3�{�J�K��T�	)�����a{��b��*��h ������|L):�ѕ�W�j���@�l~�a3(�QP-e�D��O#N�]��hA�\dZ���q�#7K��.e*(O�1�k��DƧ�+-%<o ��kS����C�}���
���E��BZ����]wFL[z)�|��z]VNԜ%���+TK~��:故��pU�~�"n��u��V3��.1�Y�W������'
�8�2FO��ۈ�|�j*����wh�Uv��X�Ƥe
V���a6p�Y��@TQ��3A��{�o *@�>��8t�>D~3���sI%.����rxH-]���~��$�4-M��q�ugY�r�]�lm$2M�STgk���Q�����m�����o��A����Zݏʚ����ޣ�6q�Z󐎹����iC���%)����'�����t`��'�H�d�-.���S���d<hi0G�~S���aq��?UR����y� N�.�*X���0�qi�g����ǔ{�ݒ����`vʖ	p/�`��i�S�zX]y�	����h$�S/���0��oXݍz[J�z��M�����u-�]R���A t���f��+ݲ�Y�dθ�T�XhӺKv~4?X���.���B��w
�$�c�����F���|�q�X��W7ӻL���D�"s8��e`:Cԍa��%<�d\߅d:���1�WG�pe��}��|v��1V��?a^V����%UD��/8�=E[����U��2>`p^,�:^�@���g�#6��"+2U!t���wM�����'=���ʹ�d'4�8�j���?�m�C(hz�^H&�l/O'c _�Vɲi�e�F ��1q�р��u1@��:a�@����������9H�BA�5�dk~�K�O��
\���j�G��l��$�����C�m�,�Q���L�w��3�ĳa}3n�d0�� T7}�U7���z�gx�&��̱��H?f�Qq~^�RG"=�i�R�fۿ����{�(��T�9�o�W�3�4�~�iq	�F����������
�h�뵘U�t��QM�zT��XgG���N�=?>`�[�t����)�C6�!؊��C�h,<`8?�9�f��#L��>L�5��kn�8���I�����c����0����Ը&�q�����"����WZ�TQ7ύ![s6ȼPg�l�c�q4'�+��dA�?cv�23�5��ʖe5�)�� c�ls�3�wπO�(��I?�1�"��F9@�%�cФ����<�5��~E��2�w��*�ѿk���ūf�6��Y��`�;jW��
Ƣ��R����S�7un�W.c�iyf�O�:���D�j�
��W39�l���CvD�p�?G�־O1W��RA�y>�v��F�ڗΐ�QH97
K:���}^����洞�}��k	|H�`�<���W���}����z�S�%ԏ���FCާU��*���Ζ�|�\Ն��jV�?mQ�&l���^4����?KvьV˕�^�UύF^�"E�o0��Ҹ�ÉM�
l���P�<�/܌�^��Hrݔ�:�s�#ѴC�"+��$U��W	�AZ!�M\=k��0���`�L����<����ji�C��TU�lhqN��-hͩ��5��� pԈ��<�����,"Ytl���+��vD��Ur7�D����)_x������0�@�+�	��)p�L����=P�o^yb�8�Ns-*�8��5�M�~���Ut�C���`{��B�T���h+���\���p��U��<��ƕRj����8��0�[�MR����e_��&Y�kj�թ�����*�ѿ�R"���&U�qe�������P�s+�)[�289�L�]9�*m�VG�rF��rM'H�֟�+v`����V���k�o��~�����R���/�Q�@�'�C�v�n<���SJ^�<���i�? aaZ9%�M�r��Mh'��)�T/��3�����S��Yu�ͱU�Lw�[�ї/s�n�m����ʓ��.�Z<+�Cا�k��vґ��c+�g�[>�0.�����ƺ�f�#&ӌ��t�� h��q����
XeF��z��፹/�}�8�=6�4�Smp巗���O�����侽�K0^ae�FP��c��6���D�W� D୴D�8f�c���K��dg5�A�H���Y�I��5l�~���m��H@�]�J9٥�@M���b$�����3��ə*b��v�^�Q/О�(���ll~+��,��ɸ8'���D*����_)���-[S��	kV_�'Y�����Jb���Ĥ����a�DW�v��x���V�e�
5*y��'��c��/z@���T �
��㝵pa>Y���g�7��c��L�k�S�>�|�x����,�?�釗r���=��6초ФM����q1�̃F=E�Rl���<�F;�Y*�~���L{��n~��0is�z7�iFa���Ō�'j�Or�j�==�t�Z26Ń�FI���9�r�_�6�ɇ���9m���J��������IR����r��;��P�Ĭ���.uʸ�r�݅�85����(	3 ��P<Ԣ*z_�~�p~�۬�_�JW��/��
қ�4�FӐ~�Y�I�uF�ٗ�|�*>3�P�6~\��Ro�w��]�%*D������Ks����o�eFO2�O�%AQ�t'm�IX�~�~��;)�Wulz�����d^��U�S�<6�y�3���\�h����|�ಈ�O��/b_f����w-x]���J��{�35�U��[���C�"��>��|aʡ�{�qצ��"�X�qE�:����(�J!TRG�l�:�ү��� �k40>Xw"�����'�܏c�%�2ٗ�jLD樮�P�ϻ�1g��*m��)���'���wS�&[ëW(���3c@hʣ~��/���>�-bZ�� ��XG�l�|Ķ���|�Vz��g�i�cap.��vI�j|縘�T�}�"���g$����(zݞ}G��Y�(`��YD_�� 5b,ީ��dil*^=+\��;{�H�nG���]j|�ͨ�C��a����@�%Sm"�t�)��V�r�{�L��l;ݘ�鑵=|/o�	!�ȚP��KD�(����g��ك�[����f���{�	��Wb��F�T:v�d_�ӿ�__ZX�:NF����)��W�c��N�Eiɷ�c]�D#L�X�R�TLe��R����I��`A��CӋ���@�Dz)�|-�����iz�����:Ũ3���n�D��&�H�Y!i��,s�VHA�i��M�R������I-晁'�����v��tj���J�u��y���N�l!��H%T?"�n��	�ө:���O��h��N�e���>Q�͌\���<�����& ��|�{[���ǁ=�!9��CJ|X���`�6p`d��l�|�PM]���<�ȧ��t��p�<FI>�N@"%�R��e�餐�6g�z�I��k�%1u�|��J���g��A>.*p\d�Pm����%���M������4N�,t��;��#�wNg=�:��e�ڙBD���tװpgK?��(��.}�o�<ɂTj=���S�s��+|��"0�����h&_10E�x&f���{ܰ4�68�:�;�PRspK��QlӐ��Xq?�i��3���(7_�|z�8�?�{�Ñ���/m���U���n�C��zT�Zt�f��+B��g�Eg(C���v�}-��	Sl�L��8�k�4\��I[�̑Y�&/WoY��J�7'�;�|�P�gЅ7G��)��&eܒ��֡��PU�A�}Ki�8���nqe��[N�@G}|�KKI�Ea;4tոt��P}k�Þ�`�g
�!���t�w5�5���bc��j�O+/��:���_�-@�e�c�"��h3Vsk6:�]�t���J�f����p�zF���Z��D��V��'G L��8�1�$
)5(�΅�3\&\���\H�m��y�y��.����U9���'<i�pi.��Қ���Y9�J&��E*�gg��b��'�}��Yh�����E�测.���^:��<k�h��2�/��K**�֊����Ki|��X�t+��u��~�:s�P��b�6�{
���Bn��Xn��(��EΥjS�V&����s�:^�e��=�"�9<�i����
L�'w��������z��x��䯢���]�*�TI-aRtW��-���M{T���;{���j2>$t B�+��zY�HE8�����^oK1d%H$2Ǔ�+l�%	t�1P��k������l*� �IOL��$p�5w����
c���!�
�k�
yC��	�Ӳ�G���Ŕ?J=5�hI3��|���s�?w��먶[�=��!�U�ek���F��fa�r/���m	��/����S�#2m�I��O�8�O�~{,�w"�� h9S5L3)�Yǁ��a�ͅ),�A2p�
��v�U[��K����w�����-���XX�[y���}A��m�X);~@-E�L���l��_H��i\)�mh!*ZH,VX
���j��H�$;��~S'�'�c����Q=�� ��Jz�D�c�*�(nUޔ��[L^��٪��0�9��r�����>���&~T���ⵃH�a�ǉ0��@&߅�P��v��E(M��������ʎ�cR6�G�!�pV+�]�N�+r�O�}�_�2"�I��C�-(� ڮ@z�,�p�d&�pa��Ö�0�+;���a�nu-�ܯ c�&���O))�ä���W4@Xs�נ�o.��N�P>�����M��A����	��f{�1��\�a�%s��\"��z�Dd�V�L?��p�܎�+ {+�=�p�MՈ�SM��#�[h(X�K@��I+��������~F>v���wX���@H���R��\=�F�6HwLJݕY��<&dZ�`W���Q�'@��I=t����'�[5��i���Q������x�'|�'�8�ۥ9�	cI.���)�8|�̓��+�qI�9pHx�[�}�����jq?z��:8�(�c�==o}_~j���Õ㍪)����S蒝�$@�ר�Atb�%�^j��Կ��ؽ�����#�tj4@�e�i��6\[��i����50̇�A��B$n������&�Y�Jr��ʣ��Z\I��>-�lͽ�z�5b­x���mp+^e�����P]`����
�����Y�p�!V-�Y��C����=S1�Hڰ���T2���z�'&,*��^L"���Q�1��앓���W�r�ΌL�1lRע�tUI�3�m�B�������CW�z󭖋�1d��`���!�rPЮ8��%�P����Ҋ�d�l��=��ҝ��ٯ'A��`��V6ҞM��緥.�EX�V��������Gg�j�..TPlF�hoi�,.���W%�P`rw��܀!���L�ˬ��6��E}�}�Д`0�=7`}�йT:h�}{T�g��_,�bA�LOPcݾ8P���`i>� ��&�d�����V��ڗ�P� fX9��k�a����r���S0����7��z[c윻�h�tV~ɑ��[J��r.�r��::j���7;z��(�� ��7ȫ
l��_����᝙�->-rV��� ��h�����ӈG������,ӻ}naE�Py�{m%��!�4lUM������w�؍��km���0#�}��jQb)�(���5g�I3	C���`�>}�g���n��r���VQ��ݔ������u,^�B�T�~#\&{���=Wu�������]������-��x����_��*X�7/uF������ϯ�G�@���n�L�j���Uo���(?�"��Q������iҏƢ������J~���_���)r����n�h�n����nPW�3DT�T���#K�;�����Xw�~}ӖsV�W���c��<�%�jx�#@ė��`'m�r|�sɢ�6�t��p�Wl5zO���_�Ƌ%N�{e�0�	�-Mї�;��W��w7��s��PX��Az�n�� ]|Z2����#�.��_��a����M퉣͐=h$�(�p��,���+��O,ЮS���'�b;V�ưgI��q襫~���_�_.�=�.�s5�㬤n�6<�6_��
�~�d��(gJ�f/0lQ�@вf�A2����E�~8�-�ܥ6Lg���\���k6`l��� Q�Kp�Du?�r�=c��=�-��.F�(4���\Ea��U$;_�;k����8b�_��<�.��==��H��</��ae�>z*�`�CstqH=��b�8���
2�e%���r'N.�b�%A� ז"�{���̀`��ժؓ���ˎ6�3"i�ڨY<=N��3���I��V���"�������x�s15�tÓ��\A²n��.�P����?X1�[�����X�ZC��dDqJ�nx�C��MSU��H
�:i�F��:>�N��q�%��f{����_8'����]Q]���6dJ6�%��F�]F��ɝ�Y��e�V�. c�
���8?�� G�C�$_.e�V��#a���|�Q6 ��|�
�fP�}��~BWh�^"����n1��2T���\�@�9!�{Q�%��/���rh�ue�f
�,��Y�)[�����(�Va�����0�2�h-=�U@\�W�25�L�[K=�D������!�vN=f\�|e��ܗ�J@'x�NN�O���Ͱ��Ȅ��6�N�>r#�;'�@�t�7�H�nC�!��`���\�?�k��"B 'z%�����b5��Ä7�]����ĉҴДDUM�䂳����y	`�N��k��	A6�"���}�4q�����|+	��z_�D��Ko���n��D���3���95�B7_|�A�c����>6��i�ȃ!����j�!�z�t��{$N.�Nq+[�y��خ�3!В,*��7����j�k��}a�mW.�����L
P2Bz/.� ĵιT.�X����W�c��N�����1[��؄��ꮰ$���0�c)s��N@�{�5	��zޅ
�E=AZ.儌�f��{f/���8%��ψ�E2�}��%�X"�lkD�/Hc���Q����6�XQa4�E��Ig��#��?ST(ћ���vTY�<�����5���/]]�R�4��0}�4[�tP':\虿[��@��Nw������ɓ��ê�	�81��z=!�>�%[15��nT�����p�s�� 7#��I�lȭ�&>���3L��ǃ�wGD菕�b�x~z'����[ǘ/���_��$�k'7\mhu'N�m�2���4�5�Y�T��.���C3�х�<� y L��n��U/'.{2���}Z$�⭜�*����4<��}e#d#����|Y�)H�Z�B���c�!.�2G���5{�J���8>E��>��a�_�G������g�4$;u�#���;FL\0�q�/����pZ�e�/�`!��>B�n�=��W��r���Fz�y�vO ��)��Mv���Hͫ6�?"f�)G-�����g�z��"�����h�<����O�۱Ҝ�Ȗ�|�L՛����>j?�*��&�Y�GZ7Ɛ+���~�x��]�PK{����?��޼�;|$s?^����$�W�H�	�S�c�޶hf�39�B�ς|�p�Dr�8���
���V�"�~��Y��u]ƌsO�v�0��ln$ePY����-~m�]�wN���ډi��O��C��E�6q�9�rV��?�
�Q��)���zbe��vz�e����.�~L�Y^����iWn:Mؕ���C;oS��=�M����9��⛥�p#���c� ��\)
�jV�=lEo��a�����Ξ��1y�Bb<1�Q��u���	�ZLk�(�ր�UPX���ݣi����4>�B�6%��b���S�m���h^N78��3j��5o� ����$=�k5�F{�!��B�]H� �Q�������B._#C�?(�P�6R��wB+0 �� �����%`q��ؿ��"+K^�q�-F���p8���@,��v���H޹�~.iC�g�NU���"V�������w��4P�󊠀��D
:ΔJ��!�+�う�Y�u��zjk�1M����)Z�^
�N����y��uz[*q��ע��&"4�Ƹ��p���Q�z��`{��=��ԝS�%`A�)<<���L��͜ʣYXA�r{!���	�".�	yX�g	���k�J��d�^_����1��:��M����n?N�C$���xi5us\�`��A�ߩT+��e3�(ow���V5���7������;���n\?�tdR�����6B�1���{qC(�r���y��v�G+��<�R߾B^q�~�­ŨC��Tmzʀ��܇l���,O��@ �E�m ڜ��z���V��B�q]�OG��Y �<Ƶ�h��g+d�GN?%aA�w��ҙ���Z�b�����F����e���-�|g���
h��;���Vk%�$�ږ�`bi �Ó.�KZ0�1�|GTw���]�ȕP�F����2���"�?���e������=ٌYm|�$��v���R�Z锘�ή?������m��������R2o��|��S:��:Uh߭��0�'T.\�܄8/�'�j���!T��y�ꕒ
���M:��nZ\$+��)rD�5���洁�jv�WFR�>��E薌�϶|��s5�FG�v��rY������[l.c��fm�b�G�=�1=_Ԋ�y��_��f���Ϙ����#��[h?��d�[\2A7�!��^ /���7}��(�9�@���3�r�\���j3�=���S�h�$��E���<g��<x6a��D.B��p���9�߻G��X&���
��]2d��T�P����~pĮ �h�9�ZLd�,�Ky�V9�}�|�Eh��>U�c�`G�:F�5��O\�~8��,��lh�g���9��������8:ʲ��uD�k
5������\
���*�i�[�\/�2 ���ah��P��Y�A��.nn������cF��]@H}�#�{��$��aWm�����x��d
���@n�E�]�(d�4���g;@Pҫ�^��%�>�䞽[%i���u���L�	o�̈(���� (�?
�	��~@�Ď�n=y��d��&���a~���@���o�Mf�Yp�o�D����n��-v��[��v���wX��N'�n��S�/����h�syW+��^<�����1��/c��7rI{=RQm^ɇneO���Ȳ��T	�G&�ѩ~?�.��d�<��.��<����Uy�S�>���
[
���SQ�D�j4L�\��F�n�3�z��y�09���X�&�o����"��Hh�6D�(�Q�S�m ��[�Kח�{��3+K~���o֢� 5�����R��%���x��,�g��IU�QK��h����Ј�����4��\3��]04)��\���f�P9�MIk��B
d��~�ºm�;�j���ìKu����9I����>��>�Xܚ����˚|A���P���~�ӷ���}�y��c�{���|�S�%j�赉�B_�E�3��\b5;��3�Z9W�n��8#�8N{B�,�3��p�o"p:I	�^�n�c�E��8�`M�j�Xe�[6'���8L�DR��X�t��E���֗�T�nE0-��q5��ך�e���o�T��p�M���F��&����;�n���E�/�����_�9�	�{��t�L yƼ8����*�q��x�s���5]�o�����C�,��"�N��E�����p�dtʛ:gr�qQgtjT��~Ś����]G�=��zC�&p�|W`���=�0;��
e��) �-V1Uk�d37����������Ϭ'��p��_��K	�{,h���cN��7����:�?��A�E���vI��3MQ-�VF�/�:�x�I�����T$GӘL�G��w��ZOoJ�X�X1W�ӷ&к[�����1䩕<��j{��e4������Kt�<��h�5C=�Hs:f�F)[�Y@���pn2$ԓ~m��R�_����+���^<Z��6&P��|%s�p�F�����]���������?D��!�@*�t�>9�Ug��)��~�>�y4�Z��i��Q���9��/%x����\˭A�<��n��l���UT�/����As�L����\�o��=5sI���H��%����7n��+�rX\�\~\a ���&�^Qw=�؊w��C��"�h��:8�Oy�m��F<,zF��B����K�N(:�q�����e��ީ������8y3�����@�"&�sf��$�@&���K��Nd#���ϐ����}�:����f�'�u����ba�hR0̯Z����%}�,Ϛ��py=e��2����K\�&(��2b��2y�p�T���C^�]���V�@�7��b�C=������-�iRS����(kԔ/-�����ȥ���]�6S��R��&�j� '�%���N��ݓ��"S��\L��Hѽ[���c*���2p��N���	��w�[������at��%�г*�T�Z�2��岥��;e,�]b"��#���)�M\�ŝ"1�B��`�;�8RFRm������Q"�Q	�P�|Kե������=��mͳ�$;<=qz����&R�t���-�����s^��1���$�%�R^��:1���O���=E�]	q��[s����y��[�\Z]���?e�� �F�E)^�\�>�ь xњG���� m*ZV�?�K`���2���l�LK�ڔ��2� ~��H�,���jد�<��
�3yC������l���"C����΁��,Y���H��욝(���	�$�-֬3�y�����L��8+&����[̫�Ss;"]��AH�n8��*u�ɞ��A���P�@�灲��狦wR�q�>���`A��B��6HZ�`��?-��#�]k�MH��ó�F�a#����fh:�:P��^�'Μ�@��"< _:Ô盀*Fן,�5,-g\�꽴u#��B�}�c���Qo���VEzT��N�H'@��/<�{yT�i�"&'q3�7�.@m�M^%&a�,�����wd��,K���q��h������O��E��n���e:S�q���\w,��� $ v��S>j����:�	���L���M�����*�����^0�S���d?�����Ee�G�,iak���4�P��g�	>��䖒.�=��4U���G�X#i��(��J(/Ɍ<˻=_�{�����I_T/���t?l&���)BB�� �4�5��p �8����I�4��W��$_fG!�3�\���L(���Dߺ9G�k׭ؿl��U��lt���ދ�&���:��0�.'��	?F�.m>���=�e�Uy-�����\#�4�������;L���̖
�.��x������C�wnG�of]d�QZ:b�9Џ*�S2u��"�\��g;;`U��·A�����]��#�læ$!5
�x�ݘ(\i%%Ӹ7PV�푣��C� j-��=�R�}��ŉU�R6�m��g��|��=֊�xH�8�s�V;����S�(L=kƘk?��Gp�%��+@�u��2�����5mYN~����[x���/��n�f&� �F'_�)�b+�~>A���|]���EK�i@���]�wȝd LJҵ!$8�֥�1/�Y���=�$�,�j{t�`�
�]����88��(1ͦ�c�l��������w�O|�
���nЁ�t;�L����=p�O]��Z2+���l���`V���Qk�����>+��9�d���&_p8�1{��G�5��x��OE���P|(��CM=:3���E��@�$�߻��%ٸ�f��k��`����������%�.*ˏ��g�3�R��%�#�rB��D��:�=�@����t��%o/c~"n�����g)��ܚ�]�o�}����L�~:�VLbC|㳺�����8�������Ib|�:��`:��ا�7~x��U^莆��`���?�F��,(M�-��g�&�N�	H�E��G�Ķ��S3�-�M(���H�٫̊}��U~��U�qǉ�$�n�,�d��/�4�fc{Z�z�x�(��N�/��*�HԿ�ӡ��e�v��T�ʮ�����jՆ����pĢ�wbch¬�$v�g�G��8�R-T��xms�ez�����l�UG����a��)o/����� �a@q&0�<�fQN$�����ĝr'f��tP��?��7&3eT�03\Y�n���~*=�1��%�}��E�����V�K1gZ��C���(d-b��k�N�O��0��le3n�Gl�g88��;�Jd�w/��	��[;�5��Kp!�t��]ŗ;T��a{��l�^�담�e��ej��H{%���m�|q����w��5�ʵ޴�~�P�)��M���p"1ɵ*!�cD$x�'�oT��!��g��xhX�V}�{�,�$9a����=�ޔ�8�Df�]�j�n�IMkm6n���4�`Ve�eb,�9t$i!=�����Z���1{�F��V��J��\p��Q�|-筙����;�|�C��`]�qg�]���{���� v���##��5�'p5K�/Kb��o�fi�=�w��yB���#h�qS��y9R�1G���m��~�D�VH��%�Fs0��A�\����k���	��_��$��,�_��dKz�\��Z����sC��A����tӠ�id���k(R^0#�����i��{U��Dx2��>(�܌1ߌ���iƇ�/��,z��U�ӵcm�*���*�	S*=�W��{W����`�&�]ʇ�+4������ov5���Q���[�i�ٰ�a�y#�ǖ�M/:�+�SF��%������2�x��\ݓa,#z�X��&��ù!�f��	7�2�ux`&��@�C`����?pp��������F�Xy����x�ًy�n�;&��eG������ֻ?�p����]��g�H]ф�?�l�J�栄Qĉ2��;�+ǡ<��n��k����;J 2��ȱM<jQ�"��t�A\R��)E�MfXʉ�)}�,�FC��M|αZi	��p\f��ihs�l��M�aEL�n��D��0e�1�a�}Z�!�Q�^���'����)����E��x��&��j���u���93W������	"�"����3�m��;�.v3M1�󥱓�}��@��d3��(�zJ�j�A}��pr��!��P���Z�����t�	K:l��n@����{�F{�k��n�WU���)v
�E�=��x�9g{k*� II� ����0L0��7�uTYJ�_�.X��K.�w)6!����վ�A�yq ���4%�������y�^c���h/����%�j��cf15�/�����	$Ŀ@��V��ތ����n�S̪,�p�/Rjw����p�hnʇ|ѡ���?�*���>]I�kZ� ���k�ӳ�S�Ÿ;ۉba��T�Ӌc��o. ��~)-����5��W��*�c�}�m�p��ٮ9.��T"����AM��ON�(Դ������wk��.QB�{�?����*�V[ܣ�c�ےpL!���~�(��f���7)�r��1V�H4⯞O��q ��_�]�cڇӚ�؂Vwǡ��&�o�'=��0*�q78u(_.�)�8���F�>�K����܂�xۿ�x�X��q��^�؃>���*��"1'��(M�b�%z���
V��`��E��d:@�0���[o���j;�7V��y	,��D�������I����H�g��N�O����R�O�)���n,�f�>:o�������e�z3�f7�U�<v|/(N=�r��}]/��:I8#�tɪ[�~h�i�;�*�}A�-$9����ge�Ʋ0iϤAy�5���O'��:LOKR�u�G˖<��Δ�#!�t��=_�;c�EKQ�4@�4�ğ�)z�MC�I�*HB�P,}����g9c�����Q�Z�C&�k�B�%)�����a�¸���)͘K�lV`�|��� �y;n�4X��V�19blz4���S���@g�oG����=8ֱ4<��N���(�ŭkLd��P�d�{\<gt�	�ޱ��!D�b:�' ($v��_	3�V�<
G�"HE��~��k�����Ѵ(�L����ab@�t��$�S~�s������ۛPW�_�Y������.�f�k[bn4��V+�[� 纑 �9�nװ����7U+ٻ|��N�A��~aBL�ڜ��xF� �v����A�}9�՜�&A�t-�Es<�Q�Hu���a��Mnڎ'~L2i���P-�����?o���$�@ ��A��;��./V:�m��U�U'��ɪY�I������|�����Z ��.��'"a;���a7�Gݷ������ğ��y�t�L� p����ܲ�*��'�E��fz�i�����oyMv��MKV$�:\�A����C*}���o3�Njm��>)�1�뿴�ac������V�|[��K�N0����0�wӲ�D�����E";��y���{���hJ��A<��o���7-ET�Q� ��ˍ�W!l�%tF۠�'e��ns���<�M=�i���au��.6+��0�E���y�]4:u~��kx�I���\FXT�E�Z���fN����.�F�|���r�!��~h�z����3	�L�u|������)�P� �1�Ƽ���N�O�j>PV��S~���+~� /��Z$�����U�[;k������h�R��Q=�I�(�~n�&��D�u
�_|�!!b�K��ehn=� �?�_��ݒm@���l��rL�D�k:0>]%���%7�f뛃�c6 F�V�ψZ���3�wp��¦3:�K&�|N���k���9�=�dh�=Nԥ_e�QD&_��x��0���D�,o8w0Lix��C�]�ˉŨ�ZL��Iw�ߗ]�<�7�Pp�x�ˤäa�(2��$z�iøG �L��L%m���.���ư��Q�.6��L��J��A�t���[Ò���g���2?�쫮��1
�'{E��u	-M<��B��ߘ=;E���^ѱ��,G������7�(�㾉?���2]&o^��/����t��3� ��M�1 ��R�$�T�l�l�Br��KLo�`�d�{z�ꕨGP.�G��z�f�^���L�[�y��,��^�%a���<D��1x����^~� y*�h���p�*5���P �]4F����{/���Cr�s/� �CDX�e[��1�W���{z��a B�or2����;P�g{��l�$��o�@+yt�ތ�+�hu++}e�ע�""U�׻�6��NE5�X��so��Ȃ��+&ꒆ��u%�NO��g���9��t6�K�"����Q�I�(���Z:P:X�N��L#�@ˀ���s����Ť�����%�.bPߒ�K7���4:�abXm��r����\�������L���!+<ǭ���(��O�}��kɀ��{�^���"���_�25�3���t�&h%��'|+�7��^e0 �A*��|%U`�]��Er��g���l�{/2� MOz��=�
�EG�8i����3���0֌��_�&D����R(��K�_��ˢmP ��ޫ%}t!k��8��I-��D����(U��9�~KzZ`*-4�ku���$
��n$��u�n����*G�-rʤ<�G��~P��<�'O7NFOe�*zZJ^��6�U[C��03P�#Izt��깄*;��Nw��Oe�l�H���.^d@�9��v�|l���s(�#�JU��������&Q���Ni֮�o'���9 7�ʭ�%'�$�.�~FV{;�$�us<TL�_;�M���^�
��̪= UM�?ٯ���na�9��ށ%zM0�q����|(ųZ.�2�ƽ�8ַ�'*�R�	�m�:�����s�VhR� �JQZ����)d��L�w=�~1:+���'A��r�ha.�Gj��4l��]9��kq(7��,�T�M�55�^$n�����L�y�@Ns�%�Y7��ȳo��,�W�����ڢ�Y�`� ����7�M�o��X�V\��E�J���̧�TZeyC��K�H�RQ�?��S�)$�E%Q*�5k��-~%:о�Μ�C��{�:#w��纙�v��=
�'���I�<���6�a,�f<0j���ڃ��z��W+�}	H�	CE��6�M�X�`�������L��,Y������uaS��̨�I�^���L��?L���a�َA9h�*A���=.�������B4�;H1#�`�H�m��#��>�z�b�x�Xm�qȅ:�1A[t��;���'�Dܚb�y��D&��e��L���ܗ��oQl�Kg[����i�6��A�Kn���y�Q��@ɟV.�@��X����-S���A8�7=t Moc�h�^E_�:��@q�	�&mI���e�V�q��0Nc�'�
�۽A�X�!gZnJ<!�*�������h�;��F��Z�Ou
\�GTD�_��Z)����7�K�\�E��3�lB���zBes�Y�m��E��G;L��?\�����1�AL�ʬ1�Ust�����P�][j�\��Pt�F&k�A��Y�����>඲e�`���5� )�]�M���A-�Oq������1�%3]�H�ެ|ǶH$�Z�=�!��[�0S�[ك{;��g��*޺���\�alm[����9�'PK��ܽ�a޽�����^�릊P��RQ{.>�QPd��$x@���脣F��!�� �zTVg]8�D���'g�+�a��KT_�S��Ώ����ҢFj��Ȇ�׳�f�T��J�Ha�����M5��3�XȨ�������K��:|�a|�x�r�ZeB��o �QJ�{�Wp6.�N���`�/� ���sT�H�PFB*4@X�B�l��-��|k� ����.��<=�ˑ���%�N�P�p�/c��j怚g��FP��],UFt�[�I�)���rR��ۄ*����n������5u1@<�%�]�}��d̑˗x_�[�xz�hq/qD�$�����Fȉ	��{�N�a��^{8�A��*��-6�w�g9��S���.$��EWG��f�>�tǇ��T{������=����6����� �Ӑ�'�_� �������9@Gr�³_]C�]��@`��@�۳K���ǖk|�p{�괰y��r�1�^/6��%�w�Z��ysx
�3��W��6���$�X��<��&�*�AN�C�E�,.��9�iR��Y���K$��v:T�A͐!j2�r>Si��?�?��%�;�?��T�^��sA��!�i9�*4��}8S�UU��b��N��K�kG�������1?U���ڀ
��(���J����c]�)eJi�@������Ր3F 	!��_>�[��b<���}��\b͟�nf��Sn�Ԝ٘�j4u@i@<s{��&�~h7�6�����-ӷ?��
ވ?�<�#K�T�䠔H�%���8�K���9(�{T�[7JH���5AM�e�w�A����X��l�����G��eh�m��8�we�L8
���$�*!{G�`�_�C���CU'2(V�&��,��)y�S	�`�u�Rd֌�/���D޷$�?��ݮ�R��/ͷ[�V�03a\��H�K%�8HX��o�S}�;��]eG�o+��Y�u�''"�Z�TH��j�aY��+����'�1�F��\��ok��$�ɽ�y��D�Ww�k5��_�e)֯�o;h�d��	&����wi@=g��aN����� ����9	~�V��� A� z[�=� Yh������Q��q��2[�X.���~g^^dAh�b�-99��)��'eħ�4�ʾ���LC�$����h�=�`i�d\��v�#r.7>��7����ǜ�&�n?Q��������;m4Gj�;�+�XS]���`�-��)�@�@����B��>�_r�k�^ �ƻ1�_ܫ�Z�YH'VI.��ؠ*4!Ӕhe���D�ϑ��s������@� ����5��/��ݽ�_tZ{vY�t��捇}�$]v���Q�p�"��n�L!�g�[ϔN[�l��Z�T�̨���EcJ#�k�c���.:쥝�d979��@�lV���͵M�nZV���q-K�a�K�r:_B��B�P����H�Rj�
'�A�������	}�#���A]�K��p�v.��/�|>�e�]h#q��H=�e!p�NM��7>�%E��q�]j-C+��`E��M\��Y#k�������3�e���6:b�gD��x=�JNh���uQ��>o\OM��������^03�\���$�#�J{�1�?}V�:�>�.���Z�GA�3?��7ر���U��pƂ��^��Ͽ���vŤ�+�|XALa�ȢM4��=�9� {@j��I/�/��C��*E9 _�G0���g
�%����)���8�!�X2���7�f�����f)��@��!AW%j�c�"��J3y�5fȕ6LB�!Da��]�(�V\�gV��/i�@� >�%�/:@�9.k}�07����Z<|8����P�~����_��7Ng OM��j;���S[&yv��_6Ȩ-d�w��+�0X#IY��cU���t�:(*���ޑ-z�B���V��b�d?�ms�̈́$�	��Ë�ʫ5u������~CJĥ�*�|}Q��ͺ��ܛ�� �QB�sT¤�4�u��]}��,ߒ�  ���v�F��c؋�$Ξܚ�P4	o�e:�C��Z]���քm����@{e���d��w���8۰�3g�ٸ߁�P��olTb�ӝ��k	ۂ��|�R
�ʜ�w�����"�8c�w������Iz�c��M�@����� %�.4�7��yi���a�Èe<tp�lȰ$��L��ǣw��,��aܕR0B���i���~��6
q��_�vYG�Y�G]���ťT6�4{�Y�|U0J���Fwr��։�����T��(���j����a��y e�e����$��)M���n�B���I�W M�$��b��1Ƹ�;���f�W9�}�s�V�l��"h�~�
c�p,�i��!��������s��$��ً��:�hϰC~nJ�I4�#j�L�����O3쫲d����z��O�Vd���,�	U��O�/i3�3� 6���c�z���1����}�V��N)I�a26�`�/ͭ.>�㇀�z,YFOr���a�AGK3�Z�ڭ��X�i�#���oH� ���%lJ�
abMf�0�ft�sJ6˩�p�	g�V6G�W��'��i����dz0/�L������*�cS�#�3n�uZ��hM( n��ω���;��:<O~vc'�{�)��T��W�vEhzJ�_c3�|V�S��L��f,q��e�e���M���������d�5*���dk	/�Њn��K$�����vĳ�K0~;���1+HN	"��B:��ۣ)��Ko�ݪ��D��j���ç�E�ef�G�? �a��QE�(,M͛��u����4"���-�qЊ�����L]�Q�Q&My�O�a���]�����hnRM�]JEsY�;�qm�f5�=��ƿu���P��(����m\ ��E��;�^�׶y���v�.��<�bq��f�e�8� �z����a�֞W��Q�m>,-s�R�#`�Ǟ�6O��8L�7x�P[uG� ��~�����of\�ʴm���su®�SV�\���x��<��9�*����dў(�nCݜ1]�ǵ��4C���i�n"�<#	�G����{w��Ix&�HfSxm���w�u�%���]��OPY��A���݇�R�?��^Q�>, ���9�ɇ�/{o.������ M:�s3��_m�k3���PpUYPz+��UdW7 ��^}jח1�U����A��͚pV/s�E'���+�]{����הx��n~�z�R�m��O"���� O�D^D�˰��&����e���n�Lm�����\��*u0���[�!��c��p�aE[�;$� 2�dLO�-�c�lS��e 
�����࿹�/t�Pn%$��o�%�x	�"GV�=/�LA��0 8Y�?̴��!�dM�ծ���R�� q�j}P�$'�IN���;��'g�_���ԏ�)�-b�|�����"��5A;zu�t]AD�9�ɀ���0��t�M)�<�**�����O?�yh����Rt.\��0��[�����ۚܨ��VY�%�m�6��V3-?���j>����v�Uwd?�H\"�U��+�xr���CֈOѺ^�!�ȟb���5�Q�$.���'Ȑ}8R��Ja�wzxk�	n�<��4i ���ƒ���B�5�J�Ir�U+�x!ʿ^�zi�Ut��څD)�3�p�t�A%zI�'Ѡ�ޟ�}�c�2L`x�PS��!�G(s>)cW�خ	a��w$��4�Y�5�H.Ќ26un*o�n��俴�@�zX�گ[g��|~<"w��۽
��N��?!
,y�<�{� �۸��@�w`7���M�A�m,bt���q��5 ��+��)���PwX�ɇ��.�#�����>E��6�k�%���+��#��g��6�� ���{��9j��r4�F�kV-��W���7�6ErL���]��>|�x��޶�Ў\a���Z`���3�`M��b��J�� �D�ފ�Z�y�t�:]�@ґ\�1)��Y�/J��~�P��XZ��\�q�0�����7�h��" t;�Z�aK,�; =�z��2�ea���e^��4�JQ���{�:=�g��=�HԈ���~}׷�B�&�y�1v���-V�l�x/LB3Ƿ�$f���>�UR}x�*�C��~&hp� B}�*��Ǡ:)�#�.5�6ӺI��g��$#|������+0 c �!sq����*�^��4��!k&�f��cPS�ӳd|�p��6??>�3w�@�ێ��j�Lv���P4�X/q�r���Xg^w���ǹ`�ĵ�
�R5#o�y�ٙ�-U�*ڮ����9��AY4G%�z<߿��3�
,\[��#S�i
!o�~kS�����z�{&ĮL���E]<�
i��w�H�����D�3�yR�<��k�F����9��R�1��d��"��)���/ȘZ,�Wq�#��n���>ٗ�ل��΄�@qs':�R��uD�5����c�������%[��Q?�0�,��f�CO� �Q��@����!ð�NV�.<��r,:�x����JgM�Gu���4~Y��{��)6�G��:oDv�$�LA���П]�Ӡ(ag����_��7J ��U�eE�?���^�O����R$3���#G�$���s�zf�*�j��}�7$�.SU���g�����򘱎[�U_�\�S��g�zv�k@���P��x.�� �ܦO]DKv�6r���6.	�s��C7�Q�OS�\Fӑ�<'����!�]�=�c���`�#xs%�JB���*�܈j���gn`{t�\O��6:-�6�����g�Г4��g�<44&J�߼���|�I<�_0P��z3����K�$�d�@p���(?_�\��ޔ�P�AΫ��>� [����*��J`�x��/g:�����q�t��,�IS��u���?�����=��ס������3;O��hs֔�>ZF���eRdcb�,��4���GwY �����E�0��}" J�.;[h�p�1���4\B*W��a.AP<��<�}1��Z�l�#=�˗忥��!;���9Uc����U����#�2޽}�� �b>g�>{���!)�\�<i�l������r]EZF�w,�L��L�fǨ�Q��BVq@)�[bU���4��-�k6��R:�����������N'�X��"|I�e���D�����a"��^����;�sLG�=�c�<��1Y�Y���nu�d_jӕN�Rv���s����P���f������s"�I݅�v���ʕ��}��DP�4��Q�#�B�%xU�j���X��L~�nF����x��U�6�tߖN�Qx�O���,�X�U����'9x)@[��j��F�=�`�����<�<����x��B{�R7>\٢��@k��++e�^� �[ �e�)`7������ՒJ`򾄦3+jJ�wG���� 0M6�~F�#(,�;���V���1�0q&z,#jy��o[Yq�����*V� ��9w}�)e� ����sy�DݘnZ7b�N��{=�Z�K$��Wg,�a<r�q���coB�tմ�:T�Act g
�Mi��-�w-�:�E>$+{?���+���TZCW\��uX���-�_��|]b�b$A��_B��$�h
c�&�[�|�� �P�Z9�N��]�T?��^'�@���q/�1'�Վ���&W|P��TO�T���)�be"tĆ�e��$�vzx4�?��+	iS�x{���nyР+$���7h�f�ey����ꉿ�u���8]�m��ǀ4��ݤ��#p4����ػ�4��M���v�^���T�\�����r?����𲲋�D!l�У���L�D=C�j��n̱��[�4�G+���O̴�G��Gra9:x;2O��'$�7��T���P<bl� ����jW��G�f���;.����AovE�I�~�"	m��ܤ����;`�s���X?4�ې'�-��^���MT0�;<� ��kS����W�a�L��Y%�j�(f�1B*8��K���C���H��9�Y�%��mq܉6�:���u�
����)�Bn7Y���	_���N1B��_�&�2�6B�RD³ �O�I�ls=�u��
�*�oE�;9#+���ho��cQS~B�qxw"k^Rt���R�W�tH����m �ְF�!�1�&���ci��J���u��(�?�-̑+�sh繒��a>� qHzE�@e��s	�ㄶL�P�@;L$%���У	�g7 =��0e���C{3z�����M��]�+z���?#�ZGPtp(X��F��@��x�N���\��@��ȟ�&�*�׬o���������Hӄ+-u�V�$�*{�P�@�*)B8���4c[)`�u��L�!�8�����S��C�-a�L	��/������PX�4������h��%K$3(~f|��M��z��hh��.��j��Ub��v�fL4��(��Y`�
~�,� �:��W���I���4^VP$w������:�"�m��?����-���%�"h��P�͊y0� #��F�:��Z<�~2)���(����{��������Ϋ,�@��j��g���tw�#��
��o���ɍ���9�mOL)�%i@ǁ�=���UG�"��|g���EM�_���Q�ɴ��]	I����vof�}��;��V�˄r��]�J!����ȎI�'ZAJ��/=>J��:>�υy<鋇XՎ��2��e���Ð���@�M@�Cf����H���|���#mX�CqDYFdZ�~4���l]e ����ˣU����bY��������Oo�F	N��5�9u+p�Z�Ж�3�Q�m�x��9�'��z@�ه�d��%֭oLB�0L�4�.lB����g)�8� $��VN MӪ�f�0�IͳB/���0`���0WtG�C�$���#�޳�-��/�U6ׅD�J� D�su���&��94�،5���*��_�O�e���P���\�xX�^d�Ғov��`�Ν��
=�a�C�?�T��-��w�6
'�<Y���$7Jܑ�1���4��w��×�q�,����7�9�ɟ-R�������ω���#|�&rp�ξ`D�$ p� `s�T��h�Ep��b���J�"�V3yRmEg�J>M�X�h��u)�+~�8ʼS��"6k񈉐��*�m0~�x�}v�	
�~e�^�Y�\i�x)�|C�o��������;��=#x*����S�	(�_��Ɲ<ݗ&猟�3S��;�2UvG��;��� ����\�zWm:��pC��i�d�(Y�}�c�qX滒^������X��pp���k�9_��`bz��R_s�J�k2���2|�@��p�VU즔$Q���1*�i��+��eʏv��Ͽ��o
Yt��*��%M�a�.��$���%�]9�d����c��������4ͼ*6��_�scl�|�t��� �4
u�@��M<�>V��\u��n�8 �k��0a�M�?��5���v1I�q���j�㧆���r���>�d ���JH7o&��Z�3��t��q?�0��������3��!L���\U�J cs�m�b���ᢇT	��]��O.4������3�\��hY�nD�B��.WO���oCvuv̦��+�zv�W@�M����>@�4��=&V]T�:$?"; �f�,��;� �w�,^��993JF�W&���Y��׻��u*^W�8]�0 %_���Ų*t��������?��G`YLW�=L���cu7g�)B���I��"U�����&ckw��ꄁ�̵Zb↙�>W\��5D#�1"�"�B Uez�<�b��?�æD����S�փl�.���D�E�߳x��J1b����k���F�N��#�,��R_��,���씜��#�ʻH\���;a�t`����	��^�ͱ�4���rn�z쨈F�kb�����B�c�Ux���LO����)��"�>�A	�<:ӳ�f� ha �ro�Q��D�s���u1z����~�C&���3�@.��߇U�sh`̵
� ��	6�R@�t����b}%%JI����nk�J�.\0� ��<v�
:���A�!޼z�ǹ;��[��*��������\���Ui��J(p[�B�|=��ͅ�fl������̙i��7GƢ�(
,BW"D׀!��T�7 �B���D��o�Å�a�Y�5�̯䇸$�. ����
2���đ+i')��疱���=z�8.("j3`Nw5ؙ��!���DZ\B<ڎ�9j���F���l�k_�ݬB�?��6�P��K�D�A�
�ݪ����IDA��Yy7��ӂ���N��'ik���v��8X<K���u,�֭�4fU����󶭚']ک�
��ů]����h�3:�3�����f��P¤�����-�G��"�HÚ�`�vṊ�$ ��>�k������H�E�@u)f=5VG6F�H�9KLr2)D~ G�o��!>-袜��~)eч���H�0�� _���J/�������J��O��,=�0~C�HI�����=w:4�U}��6����0�Wru0��X1b3�
�7���u���C+D��q����\m�	���n�}��liV6n�h���]���yv���Dʏ���w�EjU����RJhq4���ws����W}�.��m�#�;s#Љ^D�]��1��x�9��S�6�c)/��j.�Uѧ�����-�6�CI8dOT������1�
���c��J����d��@h�.|$ :��1eڅ���?�����n�t�d����!`+�?���Q."g}��Ѱ�����{�͔/h�@�1C��}'���,[�<ή��h	k���c�+)3� |Q@��oC3���]nX��2t>5h-V��>���W�b\ya=�P:�>�On1��]��.�m+[��3�K�Z��q��@1��ʳ������(�j,�/T`��g��h��,��ֹ�"�N���ZF�Mߔw1x�	��(�>�֙�52w��%>B
�;��=� G�X�NsG<�x{���V���a45��{�w�zuC�3su�Ev���l�:Pv���)�*��{""�+�_eI6F��V��9�X�ۇ+%�fX&6�X�4�.)�K-�P���Xc��>ĥ�^���Eq��Ujz}�z�o��x� f��O��r�B�eSƱ���}5�ۻfC��/���y� �t!Nm��;I�Yx������P^��!qC`X@�B�%�a�1,�'��C��ߚVu�O|�2qz9���@�w�.�U�#��M-�����lS�SѴ���	�~6�TM�i� �Bz�r8�Rq�!�S],���Ҵ���q"֎w/��m?x�����-�܋Ӑ����4��	�a������u�a�н�į0K���ʓ�zsps*M,��M���`�����X�ɔ-j3A�����q<Ҋ�#H
_T����~yt�Ӈ�k�EY�}��ki��A�@��ćOcR.�/. KhXɖv��X��A>Qv]��&��=�����n��M��B^�����JX��zKUf9��Ptu^oGlL��~�
������P$4h4}cjp�uڠ��4�L���8cĦ�Q��:-�l��^q��|j���	�5�ٗ=�p�ǿ&x�����1m����K��K6D�d�l�|p�,}�'T���j0.�uM?�j���*l�Yu���H����iku�+��Y�m�D�9PC��>#�#��W��,�J��-l�Aٹk"I!�/(sFw����W6]����U�����9�f�F-���0�����i���2݀�0�Q�.��)�<��؁^ 	��s�Fqw;��U�߱0���,G���Q�e([ ��2����[G��i��"�� �;B�I)���S%���Sh_��dW�NRhw�l��f�Y2�e���m�.鳹4V^�P�h�H����g�`�ø6��Z3�$����F7R�N�vr�ɣ7���T-Ғ;2�v_��Le���8][&��1]\0�-M�_�E:P�TF�N<�r+
�D1����ץ���1�O(�8���&���Ք�='�6-d5�/���ic�IŇ�AZh��r�	����{�G�h��	�5�C��`���<���AT3�+:�ף�w�q��ƅ֯�輛z�L��j԰��h&�ܘ����Oc[�f��_wg9
�@��dyV�yM|� ��Z��ᄅ��v�>�A�k�2C
j����e�կs�S�˰�Oan�C�&2���-���j
��;J8�|Km�>��9����� �aIui��r����o�i��:h���V��nH�Z��0I��	ޤ��'M��t7��z���L���?��=]Y�ST�|8�P��Қ�.�9�Gڦ�$��r1T��o^��	߽ϒ�c����B�%A���:�:?��ճ�Z�w@U�`]%D��ϋl�`���$l���p >������7:4B�ӜbԸ9�w'�[]�~����m�`�`G�dk�(���~/�SU� ��珱�M�a������(8{#���q��+��	.���R��S|�o�ZB^�=ʉ��:���c#4���ؤ3�6�HU6��0�����o�D�?�>�	ɠ�v�,���\G�w�D�z��0�ί�����ųDg�a�@K�U�,a���uN��)�lb�c���P�(N9�ro_N>�:������>¹� ������r���tx�'�֮6̯��U��hgzn�N��צ���Ɉγ2��8'�>��r6N��;[F�]Ue=�ڵ��W�ߖ���8C��T?�oU�0�Q"`ҒMgзdl0��+��+:��A�ă��[�I� +zI�e�v���U*�GH2᥮���C{k�Ħ|�'����5���A��٦���Ќ���7���%�ǭ�b0.'W{�L��8�H��d�Q�TQ�[����3c�->�N7��
�I+k,� �Vwt�4�W��/��籅cel����ߧz��d�dQC�U��$�S�`��w���kĞNШ�cyuI}�֧#a���մ
'Rl��e���F�y��~��ʵ�X��:�.�W��Z�O�[�����K����lE�:p6%�HP*��ȓ�dV�����d�?�/�~��y���{I՗���B��Xw x���B�{��z���#�K���ΰ�N�w9�[TM�r�L���� o������Mk3Zf�}�v��=N���ݖ*�>�[��EV?8���)�cﾧ�u�\n�BL��oX����p�p9$���R��zz��E��{�T���x$P���(i�Ko['N�P�}Awcҝ�5���@��)@�>h�9_.�%�N�U'r%�B�_��v���1u�ݍÎzI-�Q�'��.`��j�Y�P"�O�c�8�S�� 55��n5�:���匇5fv��ҭI��� ~ɑ>��%lp:���eM�ti���J��#=�I-�)����ӯ�zwS��j�i����B�\D��V@���"�����EA�$Pe\6��3�X���e��5�D�f�����������"#W�_���y�A߸����j�c�F,EBG{8U�)'���\��Gg�V��+jM'�z�����♄�[m	�#��S��f=N�����<���Vv���pQc�!5e�i�7�'���u���j���(�dRf��$޼Ԇ����	^�Ό�4S@)c��A�>T�iZd?�N+>$;?-t���	@9w��	�}�O�:����*c����[WE�,��N��̓v�ZW��2�H�`WW]7���NI�� ��}I��8�j��?�Ty8e���X����h>�� �L�ET�~����s�+��H�;�E>$�Z��(~��-R]�ی�Q��SF�����6+m���P��h��i �=�?o۷i�ĝ����^P�$$�n�:z��vz\�p4(,�f���!��U6uX+"����F��c��츕���v��xA��n��7��g��T��`�ہ�����P���վ�$�^��Q ��-�6��'Z���B�+�����`Xu�T�����
L�l���pn&�\W�_C�=�~e���X���i�����a������#�nC��T
#lη2��wmw�	GEɫʵ�t�b�,�On�X�M)Rucꚟp�]4���&|S6���935����B������-��Eފ*LN���]��A��l�B��י�3*,KK
��g��l���ҫV�<g$�踤����ː�3�ZQ���=��Q���m��u�*ZmrE��K�@A6�٬��B���_`�f��# I�7�L�s��n;��Catv:���nI���K��y��Z���� ���V$5[��ZZawp`��\��h���\@��@�Bn�������:�D�ڊ�(��>厵�/P��4"�Ca��R� /�i<.^�ByЮOrb�X"��ӥ�L)+��2^Ä�0ʨ#���2�^!N;�?� �ӗ�3�#aKVS?ۀ����St"�`��IU�W^��:�k�T?����Ƞ^��dP���9�?��c�?/f$� �߹�.@���Fdm���{ٳ��e�!@�pI��KqI{�*�B�>B��i�e�o����Q�=].����ԜGZR��M��: �Eg��$�@V|�,Ct�젗���G��Q�>/3
����������bE.��m:=eqP�j!��S'�S{�2]���b��D���������T��D�π�ףC�K�Omw|8��"�������l�E>� ���L�� }���Dg�[;?�� ���qg;L�U�������q,���9Q�H&	G�T�5z���]���k���[]����]�l�
,��v�^��y
�d8��݊g ��#ouj��Za�L7�bWR9�f珹��VY'���%���~��>r��.�������r��ɭ�l8u��r��yK�G&6��!w�{�jD�r�����!R�]V���-����g��V�-E�yC�'_ӈ+BK�/���_� $��'~�`���d���~5��5���+G��-KM&̦m���=��a|��� �gj�0Rm�xx~�|��\�!�?W^�� IT'uڜ��Իtp��oo觷��t
c��Y�U�k��i������+���0���.�a�=�6�͂�9]��ׁ/~ys�f�}���b�o�:k���8ۡ5��8v5� l�J�#U���jB�	���(4�+��IGh�h�v���h�i�G��P5#�����h|����ԣ<=���@�0�:���h���tL�`%`���dϔj�7uQzM����7O߅�ˊ@R7�=�?ի�&�>�2ʉ�>�^��n����Ov`D1�+|�rf6�6��?�P��۩ۏ6OS{�$� �^�����z	sq��3�Q�)wD.ts.���)gI����Р�����x���2�
����I��;%��x�.��)��Ǝ�����:PД����R�� ��)~�T�W���F�ѾG����@�o�a���%����O�4X�1@�`�[{��b��h��~����U�$6����n�2�m���r4�
ܒ��B�c�Gd6_ W�݁�v�������x�2�K���[��H��s|*��#5�i�W �RS'��S�d�z����δ+I޿�*6�a��5	�,:�;K
I���Gz�j�Vʍ ��h�hD���\1�\��"Pl)A_��D��_�Yl��?z�G�j�rը](�=�{���2�Y/���9ң�u��\�����K�vAqqi�݇���~��a��ݴ���?�|P��]�"�H�sk�
O���O�z��YҒ���=�i���-c���&��qg&��������X&�+@_��[���|�g��<oi~�r��Z��rC;)�㜃1H�^6+<~+��p��$������ I����i���S�T�e���{��x�b���J�ë9�n���PG$&����p2?�y���|f����F�l���g�WVrt��z��qЃ�Q@�`�j�U�c���us��+iB�ډGB����m������Ί�����b�p8�-`4���`-]m?Y.�����a�͍���	������l��Rl�Zx_��U��F<8��k�}�4��j����3��rW&4ܫD-�z/ՔLА�Ѕ�+��ѥ��}(����@R���#�U
m�;�ظ7*���ӧ��0kѨ��Ε/D���n~���9��y�Z�d(��}��~���=un����=�^g������;��_H����CS��&d��wW�*��}U�ƒc���]uR��N[�քt��	�!�<P�ǫ�KȤ�&!@����%̃�>~T�و2�8>���{���](���{{L��/k�'��8��!�q��
�����2��N��Wqg3�ғ
��=��]��l^�U��9��O���s�"~}��
��g���j°n�5/GJ�����T�-�H���!T]&_�B���;�d�_	 D����2��0�ެ U����B��OWl�!T�;���@�y���T��Gрe��BtX���8��PU\�����^�� ��͢a06��B�g���L)�Y�(��C�=�|�ITʹ��NS>� �aQ Gde"U}�>�:�,��/�R�ۦ�ͳ��Ɵ�Rg$�����)���Y����s\c�wr���0�HѥZ��GQy%'$i�t�S�PS��?��2��v����8qRrH�.Y���k��o���%0�k]�<src����}9e5�����͝Lkf"�AV�
c�E ठH��2E���hl����{�YmT��qI*z���f�M�ybT3W%h�]�!^���SmG��z��X��m�
0�<���8�u��+Jt�[�UcO��V��0b����;(�&y
q�����ph��E�f��c� m`0Tq��d��"~P���UH�*�x����ً�����v���P��(��0/��Ǩ�ɓM���0J�l��,Ј}�y��:_+�o����~k���>~��S7G����A��~`A�%��]�N�i���'����W��^��σ�VP��!0�ߎ$�7,���g�냨� K;?��G*c�E=�'3�����F}q>K>9|��q]�2A�aC8^	4^��hA	ۆbU���PE���#of#F1�B�,3c�y��r����
w��$��:�m�I��*�9"Yyߚ���xQ��}0���BҌ9�{�E��]����(*�^!�ř<�Qo�~(�y09`7��ۦ��3X�m�̘+n�������T"M {_?�'��MK�,�/B��������E5\-�{��'*�S5��JH߇Í𞻔d�3����a@��3�J���v��q8��`D���@<ϊɒa�x.���+m�^ą�)_����ut.�SAs�ZÓ>ˮ5���C	�b�QF��{����{{�^���}D�X�eGemD��(�"v_Ӆ�$���b����a.7A��²��"�f�ЌD����tf��W9�_����5����I���u���(�A�B\�2;e��[Í�|l-/d_��,��l����+�	+5[푽\+	 7���h��&���P.�{�_w����E�y�Otnd�BnJ�Ou�d�gb;��*�~3N]��P&%[R֐80��O� 2�M��zNŵ�c��JT=[���ˏ����^ �Y�P���?���&�L�a�{�{�ly����Ep��g>o�PQxT��2�8�(=����(2`~C0�F7��dt�Ro�i�
:~������~�����:쳪^LL�=\�����`�v���T2fG�އ%TuJ�>���8��N��phW�^�c%����WR�`D�_��q�T��-?��>Յ�Vf*�է>f��b�B�e�A-<�'*���"���J��d����cv6S �P�("��Q�4NC`vL]z��_�%�vE���38S���毡piP��gN.~6ӊ��9�
�l�5�,�SRJ=`�l	5�*h���E�x%НY��oF��ߧ;�΄)�Oދ�N�v���"�=�y������Y�4%S���K��$�N\���	�'���y ����OkrT���z�vD�X�^W-��?�^q��)�� <��w��|��h'���$�[^����f=��j���o!�����Kʙ����B����}��M(}3���9��hFM����8�͕v�ʐ`PiSs�J(|>@ �;(F;���V5,��v)c��;pj��mTr�)"C�^�~-����>�~G��%�o�h@�(ȕ(Ӏ��CT�����-�f������Ì)��N̷oߤ�.���� �j��+7Ã�Z��L�٫_�G�n��6�?j�#��������g��Q���Q��n����俌\"�m�{�Az|p��p`|%�W�f��C��R�V�ƨ�N���`66 �D��{��E�C�(���BrYVR�J�{���s	?�=���+>WEL8�1����&n�R)A�b�N�Fp��	�a�M8�D6QD���P�DD�j���,�}�����7���an�k�;d� ��z���W�[򧫰�95i�(γ�6�+mS�m���5i���w
;SU���=Nǋ�D����$u��T�Af�A�)?�Ɖ3.���l������5����=����򌇏�}/ֶ���t:Ί��5l��\o�3���߮}蚲�Z�iH�O0���<�`��n@�����&�~����9�P�/@t.ɰ�����R�\iM�uhbU�ˋ_�9hr�)���4�f�t"��f��o��Ng;RR��<6=_��b��b��6��X=R+�H�Sq~�2��>�4��� �!����#V��Nz�V��%��*]������P���x�I�h���vT��o(�²��Ȓ��i�M
-��@�z;�:W/����C�<��SSL3<���L�3֌'Cچ�"�	r�
�V���{�t#㖃t���keEФ*�*�'�I�*+Y�'f�۲p���j[k��oB�	�~0O��ʏ��'�K�R��uIص����z�E�+�(~��qi�+��x�ML��';���H��q��l�/1�ҲT�s�4�����{k��H���<g%c�7�{�LSk���4',�<�. H���<��\t��߇���bX�M��YE]�r{��*��� pws�K #~s 4 :�췏�VԪ(�Xu�`>
��BNc��og�q�ِ,4��3��1��q�ɕo�������&pw�ȯ;��,��͝���W���k1}���T?4b,��k}�#b潪}M����'����*�.�u�RnV�˩*&N��o�����������BƤ�n���+����M9����.<W�?�h��o������0?�ħ�P��
��I��M�Ȋ�����}� e>SX�S�&�yVB�Ǳ��*��<�ěߣn��[�8��6m�]���.���h��1��"�')o�́7��^�G߫FIw/���m��b�>D�z�ԋ��4�����F���|R9`���hk>@:��V�~K�d#k��m�>�Ş#��NU��kͲ�w^A�1��W�Z�ɏm�S����IЩ��,������^RP5?����;��v	n����ٺ�ݴ�v�˛e1�,��}m�`n��#�,���o�D���0��+��K9��2YB:>{���&K��I�f��BrYQY}��2O��i"�9݌�/S�_h=���7�	݂&�wdI�Z�`�j1b�dԦ����r�*�g�_7?�X.W�6hd<��!�?8X��� ��9�BT�`�o���GV8*�as�֩/�ӡhk�
*,{�� �)�Pc*B��2��u6t��HDi��n��N �-gUHp,��*�^A/� �}�+�=�'�34-�T��OF���	����i��jw?������CG-u��}"Q/<U�y�t�((�~M�A�@�j�����'�5!��8�N[���y�#޼�)<)p	��`2r���'����뙥�Gb�n�x�^◠���w����wr	��5�"ߚ2	�K�� �K>���.A��Dy�n����p�sJb���v����.*ҏF�"�y��P�[W8�8",�x����w5gi��	�%jH��p)�]�>�^��tX?܀�V�4��Ζ���L���e'�7�&���9�@[� G��I�M������g؞,����qM9�����)m;Q���O<�z�G�����P'\���ilx)�T�U�r������ҥ�r����W�j���ߦ*�O�rK�o�'�Y�q=Ǚ$���~���ncE��-�%$����m�3�n�<o��T��P�C���6W�	�*�F��)v\���`1��V����u�G_�Er�5���7<3�n8 f�L#(>�u�|Z%��R�Oښ� ��Q:�ꛙg5��y���]@Cj �r7v��V�T>���Q�Q����s�X��a��RP
�#�=*I(��|C�Q��*��y��[F�@�{*L�^��)m�H��c��o�!�8�w�2�Lѽ�������g�]�yxl��~���5�=j�����pn�6�E.�MT����A��w�Pz6�����A@P9�)(Zr�t�	�1���'V��5FEP�:/�>3�h��*����Hm)��o!������qB��J������$CSCl^tW;�q��U�����/�E�A���Ȅk@�?@��Io&Ĉ�� ��u���*b?k�`��Nsb22Gߢ���V$)�
Q|&�xD�ꯛ�`fK�Qm�q)�8����
K�X�"���[4u��� DY"�W~|�0wXͤ>f;��g1�ì;Oq2Xק���;}�,�����`�#�=��|����[��Cw���!~��<����[��AW�A$#�L�;Z]�9[�����}5�������	�>�2�C�Pd-�Y��"˟F�/�<��
�&M*�fU��{)mG��,'�l��W�m,U;�q�n�w�.�י�Ys�&'5cͺ?�����V�D��ق��v���nj����-i���<�Q &,U|�'
7�y_U���PM�+�|�5XhȢ%o��<��ⶽ�!����`��'T�.����/	ɦ8��*�����+17�>���Q9���V|:���eK�Y/=/�9/��Z3'��s�^���(��#��M5��� ;e�����X�����X�٩����f!A`Q�cR�=��j[�b�nQ�k��`dc�zM4b~y�"Eꈼ���^g��==��xQ��n��܁,��&���L��6�f�q�C��_]6�@@����X��<G��>��ۈ_�_�
�����;���@���ﴦr�*���W	-��G�w�U�>?�}�"�4��>'z��9 1�h�:�n�=��C|�v����;�m��uOF���3�u����]���+Yp<f;-Ϟ�R(�St!M�	�,��O�{*B7HT-��/cogn���2p���>�z�VHh��=�D-�j�J���\փ8�1�e����P'(���-�u��H�mb��~{��a��L��T^�;�F ��.�i�c�]�^�ў���(��JUf.���ǆ$=�b�,=��M��n��}��0�P�Φ�	�@,��h �ft&&(L=���qI-1j����Tq�p��b�?�xE�·���ݼ����7�3����PO���,$�[19x��~/K/�Q �s-tm�r�]�,^��=X���A��as���܆�����IsO����������q� ��S}@���������a��QI&�[D\��$eT����S�Dp�8�k���o��QU"������g�!�H��Ǥ�;�X!���8Q\�|���i�C�;8i�bѓ�Z?xU�'}���|!U|'!�@ a^���_F�'yn��Q��tح�@�,aNQ�5��g��S	Z����6��!����v`w�ˎ?��`�����l9��]�<X��ź��s#A�f�L0ð�Iૡ�c��#���̧�Q�O]1�k=W�O�]g	��*�}��ǚ��ᓚl������n��"�P@ϋ���g�1~���ꂈF�˕?�|3��r��y��0�&A!���v�̫��4��Or���!����Ͳ1�r��oi��X^������uMO�Xֹ7h˟�F�5��V�'���^��lu����K[�!�hP�W*��>G���:�����P��o@�#�זg�v�:����*������J����m�z�+�<�z��.�D��^F4��1U��p�t����3�z0w���{��G�#����+�Vo�o�u0�OHl�/݂���C8���}>�wfǬ�rM�5��Uϻ��h]���E�AR|��^l��37�Ѝ4"��T"��;<�`��V/"a>��r����ڪco�׈l(v~d��� �c�Ȃ+I	���E�'UG"~2;��+�ltt�D�F�if}.S`�n��dY5}��������I���w^E[q�C��&��Bj`U�q֊��I�~z��/�C�M|�������e�-k-reW�j����Ux3��}M|ߚm��ʘHޒ�!�ͬ|����T��4��jd���'�F}�P�Z}ϥ&�Z���g����'�K�@P��Xh(�Ĵ.�4/�F�oO� �|a���G
�Wh-U^�[_�u������lc�����\(�����G��f��S��@��o{Tr�� p��g��s��P���3�D���y��w�(�E��`R!�]�x���r��a���E�!�IR�����p�1Bx�&�r<J�J!-�u���.:��J�����u��B�1b��}`��鞩	�L�6���q�E�Z�t�J�<��;��p���i��v(��1Ni����vz�W ��5T�'�vK�Sd*��j�]2��G�!geRAo{뺟ڜU���6����"��u__�e�1-`��E!!ڟ T7v
���D>�}R��fy��"�(��Ǿ�s᠃�}r	=��:Շ�i�+Q��0��ŝ�er��Uy.u�%���:��o׫�ۭ-QD�0����4@#�n1,N�����*�ӡ7���������|��B~���uĦ=lA��3���MX۩B7�R��0V������D�;p'B�"�P��������*OMd�qIP~�c�1�����:Ɓ�T7�`/l󿚳�.7���hb����\��+,C��Q�Fh��)�������T.=!�h'!x�5�E.'�0�#Q��ІR0�w4t�&�����,���
������.�]�l�Px����C��!)���dB!į�9�F"y^n��3�H��W�ƞ �H��`�:�5����:���\��FS�@.��%��v����5� �D���ŵ�4v[��n��V��Gt�w7Nɳ<	�A:��b>��sxj��4�{V�C�nR4M��͉y]+�*�C@����L��5坘Ű�T,�p	������/.x�QZ{�`�7U���j����\I\�r����`U�����9o4was�ޖzc��KT�OG;�o�8WϜX�(�n����椋��g���n ʹ�3˂M;��%��ުR��Z0l�m[��X��뇻R�~�*v���H�2���~���#�7�8�q����1Ƿ�~��Ϊ2�wwEu���D���Õ��eq��G5Ӓ����,�|�4���ƯY\(R���k�F�QB��Xg��������8���N�bI��Eg��M�(wV_���nٽO<E%;�M�h��Be�2��bR��;I��>�y`l�d�܃��4g���Nx�Zb�;���2�
д�LM�[L�Xf���d��ÃøK
_��Z�-�1��m�����:S2��^Z�'�j����X���MEv`�SF�Π
4"��̓�V���O�}'!g�����n���?�8imW
�n���&y�<���7��JL���׬�	Bb�eX��Ag����� R��L�$6�'zBc�6�6Z?h�vw_�_QH�5�}�+W*���%طq���זv1-���b%�O�f�!��V�A.{��o��Q�K��S��Rῤ����a�z]6 _�y�a� �X���>(1��*�J��?����8*|V�<)g���u�[QL�HhϬԸ��M��s1¬t��5똛Mf7�  ��dId��+3�0�!(T({����`t	�y��@8��K�|c��š���C���x!������h��ޡ&_�,/��XP��=0;�,�?L�osC��d�qX�ƀHe�@N˒'d׉�2�c���A���+{U�k��svI�}n�#��`ϴ3�y~��C�H6�ѧ	�=&��~�����v~�`[/��鄭�&EZ����=��8�ψ�'�O[�N�볙u�6b*`�B�B\�gR����~��s;P)n���䑏k�8�(��!y�=f���&�.*z���I���[I�%� �((���&O���ۂ���79@��U��9��ů�	�)����#�!�ۣ��l��G��.�r'�ٚ`��V-{�̯�wGB$�q�[�k�E��Px�'	��c�ջi5�`��%����#)��R���L����$erY@��6��aO2T���v9�JkkFBc�Ma�lp���|�_�̳>�)�������#i"9�Y�[X��`ɒJ����E���w��V���eS9�d�3�߃��V���C�]�zg�G�������Rl>��ȑT�#\�}O?��/&�4@A��V	��n����4	�.�~ҫ��������lK�=M�o�=��&��K����X_�ϟtX,�z4�q�b:$`��@���BI���L��m�7��R���y5oaM;_���V�Xƛ�1elx����o�-����oi.*�g墠��0�V��k�WXF�U���X2D�z������/��J��mm��4��l\�֠�DC��jI���,?�eu���x�d8�_�iH�3Z>��;�i욍�rs���i�6w�t���T�;���35��:�k�h�i�A�pϛ]�Q�ۘy��_l�ð���9W��w��� ���# �#�f�������1�d�[7w8��]���ȧ0�&W���@�����<6u���s����7Ċ�yk�w��Dy�/ab� �>���C�c<,\
��3!I�o�d�!Z߾F;��aE\�봄 ˪��|�k9U-s򍦒�&�omG.�T���F�T��}50չ��5`����,7k��L:�&��y�PO����M�>�V�ȴa��%9��������5<�{n{����?Z8�r���P��ԙ��N�����
�v��o��s��X(҇9~Qfs�f�W�z�L�J�V~lΧ'��"����6��x��� Y���^����0B���C��r��W�L=G�xV���"�Zj���N[2`��<E�����R���� �E}�C������BVӼ�,��:6��쁀���Ց�4���~=4%?�*Sen'��p�J���zl���U�U�DF�H�'��W�j��{�������}���{�P��WƏ�*8���;;w��b�o7���&�u+��u��;������(ֆ����UZ�5�>�`wLs���9�"�  ��Yn��D[�h�!Lp�Қ�s�d��)���'�%+4�B��*��R�#��^+����HH�z����E{g焇�-�xe�sCv.u�i_�vh�k�l��q+'�ǃM_�Є��o<���n��]B���YS�@ZU�o�i;�MD5M����D�/��h-�m�������0,r5�Y��[�|���t��W�R�ֺ��5��(ϲl��%9��m��]��SPUۄw-���MY���{�<�@bN�� M/��ê���Zs�:8�%�bʽ���G�ף�+1��і���Q>���X!��N�x����#�7��'���J�,�O�M�sJKj�[�+�B�<O�=i�T޳�ߝ.Q	��[�0$"�D���Τ��4��!�F��3�o��鎑�� �/����#�@�7v��Ͻ/�Z*���ozt�,����(�ѧ-�q��%�7��.H쫐a�>ݕ~��Mnc���.h�h:�"'"�?ȕӶ�g�,�������z�<?��2w����q��i��j;���\}��yG�#~���nZ�n0��������D�Y���(m�(�lR+ǋy�E=5�; #h�.��ꨊ��0���$�;i� �M����cW�e�0�ڠ��~�q//p���S�P�(>F�~cy!3��p*1ޙ�k��Gh<b �Z�I��h7H��7Ui��Έ��D��㫷��&7�#^/��c�zguZ����$&�Z*@a���hI4��8,u]��ĸbj�xΚ[M@L͔�V\*��Hy	Cub)�e��@�\�ܟ�3O���c
ӱT�K�k2�B����� �f�5�^�}�3�MS��g)�o5���	��xS-�R�e�fMH�9`�������W(�[�ڞT��&��bS�a!����O�^��N�f��*`S���x�J�s8��C}��_���V�!S������l��EȌT���E���X��bl�&��n�9��?�l22���'����iFS)哖�����c��W��� /h�h��G4[-�,?x�����N�*��l�f�7/����:q��C�X.p��JŮ���ܪ����D#a��7��3!m�mj��x�h¢��O�W;�ǝ�,�`O�LW$)n�
����g�+��y�� i(��9�W�;ψ�衟|>�G�'�&�����Lϟ�}o���9`Ga�g�,����1<�Հj��E��a�� >k��)�a��RRw��LYaR\U�P��2ec�]ȧL �@��d׵�*�d�p�Ǝ��Q�c{�$^ĝ�L��T7���S�����Cy�>��
Y�E�1��!���`�~�M-���b��!����%rz%n�8%q��mR��ya\���Nޥ�:�R��>�����S�r2JFI�M()Fۚ/�B� TX���=<��TD{\e��%�Gkq-C�'�_U��l'̴ke�h����5s�<B�R��Jߤ���Uä��!O��b�.�"�c�ց}bx�!)�T΅f*��}�š@6�|zh�VJ��4;4>�F�o#�"�����%T��0\� ���wk	�C�\��bֻ�w�h�!�T�gwكV3tW�H��|�86�k��_Z�w$CW1���8��ĥ�0RĢ�0��{��b�5�yO�Uǈu8�=ٛ@�y7�7��|-Y�o������>��+�w ��"�a�ّ߰���y��<�\k^��q��iGU��N|�VOB��u�6U�oÀ�w�� �2^�U��牬�r��A��G�?�J����׉Fe�6e�x

[�S?ŵl)/x��|��0�������+�{���r�S]l��D��^�H���7�,�w���m�
3&q\+�y�����L�:#�Zw��?Ӊrz�f:�z�p,g�$����v��$����h���	�_��T#kj���Y��%=�(�Q�j�C#ߴ��w-x�<2S�9������{�>W�})Xc�.|�� �}O����ehI��i�/R�.�u<�����9ݤ�Aح�y��&��+��,�ҫC��j"��fW]�G�h��	~����oܘN`�����u��'f�H�a6�aT���M�%�����oP����Z����E��%Q�p��c������n]1a�Ii���I`�i�vfq�`/:n��k�I�.�{km!띥m�� �cQ0IKE����p�3���E���.h� ����g�Tj<M�:W���(+�Y��㿱��F}z
��N'�*� �+�T�{����V(�Q���P��=`��A"?+�^�2{�e��v*����1��(���[��k��ÓPr��Z{���O��[ܔ�s�?F�	M�u���X��#F������nHY.�Fw;��f^�Q4��?	��#��v�>r��?C�^ř^�����e���+��_��0m
r��@M��#�Ծ���X�,!�5H�.R�����\h�#��H��ؼ$_�{?�
���mݭ_M�TϺ�����TDL��S��,�܃�����s�� ĕ�6�c/�ZT�(�'
'
6`���= x�r��\����,��٨M�X��p���*�')��0X����&L�n��Ϊ�B�e6e�FN�O��y��MП~X��I:,��∨�(����Ob\l̓'nc%�WE��ӺY��1Q{�4a��$G\�paͥ�+9���k�C��*"%P5/��l��[�Ԗ�u��2��׺4{n�6c����L�r�؃;�p�~Yh%'�������#Pk|#r�k��n������q�B��*�]�_�8h�I#��hx&��R5k|xE��
��1W��Xb���x4s���)����q�\,���}���	��H�==�`��"Ӧ�1�ɨ�
�Ti�j/̧]��L�_ɾ����w�ہ;�LF����m�j�.��5�'�7o[ğ��Z�
Q��w��L>	S���b5��㗦Pw43y���xd̯��v&қ��΋���+�y���|\���j���8�^�h��kQ��X�;�VnE�yhg�.��k*���;zt��HU@/Ȅ�K�&���ZY�ha�^��Z�G�h]U�֨�ݎ��t�0}����k��Pi�}�p{��1*?����|V�:�HB������pEI���}���F�j���jr����щ�h�6r��ï_�+т�L��Ӷ�}���|��)��I�����Q
x��q�ҽ¯<"Ysyu6�,�:�H�,?@�Z7�i`l��C&R�,�H������2���0x�8=Q{�m���I��I�q�=�ν�qsɞF��X�d'�V��|Mw��Gx6Y#(�[m[=�y^A(�K�o�Y��Y���6mw��U�����*�Ee(��Ŀ�P�B�u�٬R�˗f���8X��$�n�p;4�7�L�""��hOJ�^w�JD�cŃ����D�q~����>0·Ϊ�@���E\9�^�븙�"E��o����m@8`_�����׃��V����U�z�C�2|!�$��Bz/�}LiZ��X��p�/����c�>�=?���L&����?`��-���,g\�u5׻\<� ��c�@Z�~���1v��I��W\rt�c�a ����I(����a�y7�U�*e���~�"|�4�q>��Y�&R4'?��pN��X����J�v���n8�H���?�xnT,!��͋eZ>U�fμ����,�x�=n/0�M�3a'[��G�X%xA�u��C.�^�-�YL�@2�}�����ɷvs�OG�#X�%��]���Z,ȏw�J�˕���\�cc܂ofC�,xi���{���$�P_������l�(��2<�"���Q|�́�H�'Ȟ�����'��'᪎����e�4� �*W>&o�sPe�	.�3[������!׊V�
Vf�.,�@� K�ϙ��~Պ��� �IDx�S���q69��\�0���LĝBQ�r���S"��P���,���m�S��	��Jn�d�Wy����u�������(S׋��sV���Ɖ![�O�Rz�Lt���Su������F���1���"���	�o���|��rTA�U>c֒�J:>�q�����p��,��u�3&gnލץ�ӛl�ہ���a���TO�dg8����F�f`�0�pՂ�:���kZ��t�6��'�r�Q9�L�xp@5���F|c�6;d�7��j.bK���F��(��>)w���қ�Fz��E�����8Q@`lIڑ"j	^
my.��U*L2��⭍Y`������B�=��OpU���"�����0i!`��*��!b�]�l�Ho���C�$!e.(�<Z#�E9�dkl+�!��v˭Ѣ�HH�(9K8s�������/Z�+�5!��G��dcWm�*8�Ċ"XQ�hh��/�: q�P�� �)�+H9�8�w�LL���x�4ƌJ�L��Yq/z�nn�B�@R*�ǖ"�@�a��bT� ���)�v�Q,���YNPGSO���l�Wd�o��KۑiI����{޻��,�_e^�����Ͻ��>we����K��g��6]���g�R�*ޤ�<�-_�����g��!#�շ�bM��F^�y�d�#(Íw��>�y�Q��#���R	�/r!u\N���@�;���&��R��\ձ�f�V@�g�2:D%����pA���M�����\��m̡���Q�%���-x�L�Ǐ�ݰ��W怜e�,)V3�>�#X깨?D�ayb��K�Q`
�l�#Pr�$�v7�	�er��9Yf��F��
�>�=8�	RJ�Tm��q�#�Y�E)���{!hXs}_�aq�n���\R��M�*���7(�J��
ڙ�M~iF�;U$��3�s[��~#â	�� �>/��T��!h3��!�!cN�C%�Z���#~_�~��k��|g�ɡ���Z�J�a�k�DS{�v#�ac,��X"�����B����&Z���t`硽t��(4w|��i��Io�=K�M�l�_��-�t$S��Y�(	��j��O�K7Օ~F�Q�+7*o%����J�Ќ�2�l7�QA����1��q��c���J����s���Ң��_���R�?Gd�v���.��FH�,�ʧ,\<D� '��C?��:2�w��������#Q����6�ٔQy�C*L$� ^`��h�p����F);��k�{$X$�e�Zɘ�y�s�Ԧ��e<���j��/;�ն0C��iL[���/��իΤ��ƴsu $_~����O�5�� �i����c�c��ۍB��Ϥ�P������&���UuS��_�ױ�s�b�f�z3��;֍h��@��ƽ�_���2���B4 3��K+�R��v��S�.�����s�Z� ٧[dZ�)F��c�,�E��h��@�@��dҐ�W<ޜl���E�ݴq�� )����^���=)���u�p��
�4�b�Si���.`�X0����N�w�%�3�u3u����D3AY�y���4�>X���d�=�~�6�����/'�l}6�(�g���f5�C�&����po��#x�=����˜�M��k�dwkE楥ۓA3�o�;�M��IP��6[S�';�&=�5�W0�7Q�{���A�"�û���f��sd�Q;2�d���G�}ۺ� N�g����vq������9��k*�s����;ѩC
��
=�1����)`��;�Gh�]�E�@��D�2�k���v����Ĭyە�c#�n��Ɲxs����=���)��ԡU���8�m���P�F#q�����S�b����ٶ���E��'EZ���|��s�l�x�Q� Ԗ�B��3�_�K��l�2Pj���홼}���P4V�]ˋ�2fRq���i0���%������Z��|����Tj ��F�V�a���Xx�,���X�b���QQ��� �jx��/�:�4��,q�r�l�N���5�^&�L'�#����u��ޛV֨�3~��V�����I���D�x��L�����|�[ȑHb�`�l ��(z"�	�l����ZUM� JD�ڏ����R�_ˎ	n$mJ �-�*�lF�Ձ�/YK�ӌKN@>Q�Gܬ�k�u|6�g�,�^������_�-/���E�*�53E>##�n
U&�<����oU7�!�k�R�G}ZI7����V�T�1\�M�yWo�N7����(xȨ���H�����9�Z09U��L�:�Y؂Q�]�E�$��eI5�	�ʥ+p��]�yMm\Z	?x���W��6_���X�URv��jt=���q?���/�%�d�~���[�A����et������-�k!�t5/���f�^V�Q(,p�|P;���d���g�9%9�r_C7��gM�w��G����.�v��҃��M��E<����L�@LP���]=]�U�M�Ϛ�[O?b�ط��DԔS@�:{�7M� Ij�LrZ��&.F��u���t�}T(��(�N�O��wK�|�(������b�}��_�� �h5�A�x7R�&�L�b�	M�`�<hQ���~}��S�_p�P�������h?��01��9�V{��̡��t�`�_�ͦ��w���+�K/^{��#�q�n�M���� ߌ(�d�X�#L�q}}���X�O_�,,��y@7R�Y��z�6���s���0�5�+���w��%S�3�v�G�a���3��PТ��w�t���g4�@��\q飻	�I7��Ceˮiq�ybq�rȲdk'�&o�mV�~����E�Q��΃mj����>8Wf�4�=��G"q\��C,���p��/l���26=]"b�˝��������`�=��r����v1��hܐ���˫r��C���`>kr����^�U��|T��n#z����jB JĨer����}H�C���2�/�H�몠�|�w�6�2��!��p!ުZ�t��nw�؎;�@Є/��%⏏�׈�r�<f@�u�~BϏW!6�3gRTCH����
��LE��A#�7�U���FW��C*�v�8��dԳ-�$�4��~��.&%dK:�Ny�wd��5XΛ��[߳�u�o�1�^����[�u��DHY1Vιz���!(e�FG@w��5�T�F�^3e������]o~��"B��+p�����9#y���?�8��kJŜ�n
�H�Ŧ��G�8 {=�>8p��D��Z	�\=��.��ӫ�w�����������4���2J|�X�'~��x5��T�d���u'͹�DP[�F8h"�#x��+;x�<c*�A��Ȼ��7dZBxf?���W9"O�SW���-8���) �ޚ��(��
3����I�D��.�32WGL_/'ۖ%�"�
+a��в[q��3����Ȉ���:|�2t(q���)l���5�%�1)U��#(-����К5�g��*�R�$0}D=����d[Z�M_B6$���Ua���az�P;P����!	����q�?�Y��<�'����Ƌ�g:Lə��g���o6�qY�}m��|�(�:������&��"48϶o Gl6�1H�DR@�>R�zy�7�,L��caU��6��I{'Zrz�1^;;]��N��Ljs�i�H��D"U���2��@1_L4�M,�İ�C�Ka��5�N+T�����v�a�`t�v�t%&;�:�/��d��}��P<d���uf��b ��[�u���S�K"q�t�O�����<5�W��	�hfʋʵN[R��.��p�U��O���ez`<�=5ر4Zǘ_��@���;�8d�)���+m��v�ϥ�ٛ�I�Ïqֶ�kK�{�z4ꪳs%�٫�$�o����?씐��%R�&�(D�ɸu<�*9" !��z�YZm�$�	W6��y!]]��hw=9R�#k=6Yв1����P���~8��-x����|��ttY���	�y$���/F	�2��? 2 �%R�z�9ED���ǚ'&Q�cR���з��ƈ��\��1�h�"|Fr�j�l�4�Ay+��@w�F-phP�����ѯ�2�P(F�i������:�J����Nʷ�>5�^���A�wYd|�������*�z�W��["�	���e1W�G�gӂTÈ�^7x'�V�V%�

���(�E1	[�)����3���2^�q��qYpw1|��a�D"�0�eb��G��FҚ|=�a.��������?���4t(L,�Gs0D��<�u@�x<i��ߨ9[��G� �6]ޱ�{MQ-���C	�#���ր"BR�}��0�a��И�l�#�|FF�4�o%5~̠��*�"�D�f��a
t!
�شI,>�����S@?j�x������F?�����"��ЃF�
F&i�P��pRT �ګ��W��dg+��Ԛ�� ?Hb�5\�r� ��('؟��� �{Z`��*��? .�T�����+�1b�s� �e�<د���~�+�[Z36m�_)RR8L&�dI-� ��QHZ��觖���4O��I�W���,ܖ&/��g� �i$A��xr	I�eOb&�O�n���A�������U�����;�HEK;[�Г�3�/Z�B��t<�����2d����4��V��Т>���e���I�m�8�_�Q�j�j�_����;��=(Q��Ӹ�e���]k�}���V�������	��v�.�;Jg�݄Jow��ߞ�#���z)-��!d�]�vUI&�gQٹ[P(�-��強H��e�'ƅL�S_��sc��H����:x~<[>������[[��z��:��LͬC(�,f�?�Q�*MFu�X�!�9�D�׎���2�l��(,���Z ��)xt�;������������>邛2��c��ّ���!g�oy��e�Y�y7?��\Ғ����{�����}d9� Wn�������;<P�)���]��<��A�L��k?mF͇�'(<QB����m������3�\���-�����R�S�y?ȰT/n��\k�6�M`�76٥*���\��-+,�2���i���GSZ� (��h��Ĳ*^&�KM�Rb��Z����ϻ+K�x��g$Y�H���k��rj��zA�7�����NI{L�O����NA3߁�=i����A�	'-ȃa�0Yϊ�Ad��M�)�%k�R���v�����t�]�P�Mz��T�]U�(�9mU>����ab��v��z[�T��b/Ե=����)C�&�!���GnY�vh}��lQS��4����9���)n����\��#�az��ȎZ������3�g��y��s�/���y�K��|�%��	��>`��洦:%��#�j�j����>z#�\�W"r��:�Y�E�4���X�1޳#���gҮB��öQjs���@�1��_�p�a�"� �P*d�$v5K����U6x��q���bI@<���#��t��q*j�2+��k�W�D|us����
b���%2��P)�"��xa��Q.O��`r j���0n|����K�Q��t*�G�Y���p��I�,C?��pv|p�ҙJ�8�i�S��+3@�\A@ I���eЩx�`ey��I�7���a�/��Ň��$KR���  k���2�4�uc��4�M=6��n{T� �����'L�s�y? k���&�vU���'�wN_��8�L1�*024ĥXR��k8nˤ'g|��
rU;*p�wS��{��I\s���}�F�Х.>�3̈́�ffF3T� X54Q��*�<�~z2]BB�Pる�5��h���(e�p�%�ao�y� !��N�e0n��)3'��=�.��}�X���A�� 61�G��x�+6ä�J��kR��$�8�ƴb�:D��]z� ��*U�;�L�C���z$�6��y󨖔ҿ�G�e^	�{��;�ҁ� 1��L��6Jo�G��Ĭ��0�����Y$O;$Obfk
r���	��ę���`�>eNf�t��sJ������l�Ǉ��Rg.EA���g��W�6�9����$p�>��p�ꌊZO�=q���_r�lt���\JQ�$�˪j����>��q�>`�� ���e9��?=Q�K��
걙����ٌ;?�W3R��a�c�L���?����Ef��Z����Uw�滴$�h�������doGg����0�ͩW��أ�g�L筅'�ϩ�3�^y ��	�y��E��Ic���uڹ�=C��f)��- ��s�Hz>�xn܉� 	e���4���BG���U���z��M<@�eڅ>�27�B�� �%%!]�e��u[���ˁ��u��Z�����d�ꄀ=��5�%4U+��|�DI'�6�2iGI���7�x�mm�E�8��Y��e5�T�������
� �}���b��5�@����
z�GԞ���R�� 
�>��b���G<�_�|��b20�� E�7	ݥ��T�w��kg��o�3v����Yڈ���í�CC'P-�8�����
��ס��]�w ���,0�($Up�E~It�L<�D�����N~%��W|S)<���&�l��ÊK|k?!R���pI`��u���U~��	nE�33UL��G�	��a����D�>5���2�6��@x�6�]��Z#b�Fm~ݣW�NI���ϗ?^�x��s���܆g|+����[5���k+�,"�_��
���
։=%�oqF�D$�N�������n��5�p$�Y�P�`:{H�]�1�W��x��k�F�R$a��k���q>��x1p��{�5�|��u!�nS�s���@3�f{������Rc�������a�p[��C�҂�R�J�y�ɇXN�`�������>�(CBT����al�᳉Z�{6�D���@.�G�u����B��Wy���tgi�� ����Q! ��_p�'��R�-��_G�)�߉�^DӖZ�̎�j�)j{u1�x�dH]_\����^����E��
�<���<�����>�H�A���X�y�)~��cy���{r��7�ƥ�[�;���dk7mx�c/�N|5q� �����RC�O�������i��W�ŭ��w*��	��u�R�Z�����aM"a������?p>GL$���h(LםV+-�A�z��9�m�S��J�vc}~B�2�� g�U��8�l�@' 6^�5l��Zf�w�!RKYh���(4�J���y[Cy�z��8b4���%v0*��t6���7��H�C������@yQ�04�M�:�F���#��{z���q9qԔ�O�9K������j���#��:8��\�&�23�˩��y���<G�.��^�����e_�~h���豯zV��k¿Ǐ��/��ڦ'!��>��i	|p���l�Ly�t��֤t&2�Q�M����ĿKM�N�߈T�좼ѻ�p'����T]de��`�.��AK9�7*`0�ZC�5H��:���ڨ��:WM�'���l�pZ�pRº��k��_Os�����s0�	e���T��@������j��H���7;m�u�@�9�P`n����������cTZ�U�x
�F�g�S�_Eе����<Ŗ{2"�����8����6��]�|�����u��⩶�h!������+��T
�~�s=�1� �P��0�����wo)k3`*Y���k�$�n'2�� ur��Ӷ�6[H(i�k��q�'km�^��ظ�A�݄�C9��
:����C�s��K������ga
B3��j�uIm�ߨ�P�ܳ�:�bì�3A}�~��'�W����F��[���9�v)���Ab���r`
��ٓ��쿷$	���K�s�WR�mA��6�0+lr�����>x���w�&�K�=J!��
�W,{�U�l� z4���RV���C�w>��0	�5-�����t�8V= |�5hj�,���I�2�"\\�N|%n����^Z�26R'����� �^FИ/q2,������?Z72�b��m��,��ɻm��kJ�י'�V�'����׍Up�Y�'��i���4�JK�d�(f|�sH��ZN{Z�8�0��Q���֐�}v9��o�l��4tz�DP���2��RQM��Iu�?���/���6`)YM��k�^�~��w9P�O�@r4�K��U;1�bE��z ���QLG��Lx��,S���BPy�Q�#���@�4u��>��{ɤoVL�tԡ9��&O�Ř�$%�.`#F��!=Q��ІݠL �Z�����2�z��,n>���a��И?h�Q�ˌ�����/�څ*�7.F���N�0���H�W�6>�����h�-�;�(Cs��N&���c�ͅzsf�kR�;���$�!}�j����(����8C*��,7�&Y�⣬&uD�c�U�t�w�_M���b4�&��t|�3@��dv�q��+t��)&��Вw�CV��� !p[�{���d�Γ�nk�ȆO��CΕ!�o��gs*�BR~yU��#��^����$����鶺�d��#Z��G����Mx�$&�X�Zy"ϼ�N%�gX���[��s�W)e��ye�c�2KT.��\��)]H��<�@���x�m	���e��+S$ҧ�#^��ݰP
R�pF�{_`k=���!]9������$of�� �S}.U�i�Sb�=a�ٯ��z��$�U?�y�kA'�@kZ�!�SO���Q�������r��~1�J�����f�t�EQsNBa�E���ܥ�φ�{q���:����l8�%̚���/�3��\kO������[��)T�)2�c�<Wq�����,�I��nJ�B7����&�-���9v�W��!�_�D����k�����6'n����"�ܣ�Kia�J/�I N����,��/t�EEc\��"����J4��������*�� ̙��Q��Q�Kf9?#�9��D�%���}g�Dt��:��nuo'�h6w�⿗�e�!ZJe}mU3�ɹ6���
 NuNG(b0�L\��V[�c�en�6 ` �7,zT�Dŵ�ԣ��a��̉o%O�׃�<^�bn�iČ��]m��@�2/شZ�@?�%K�e�L�ӫ�[b���^M��Z������̉�����y��mT�e�Y��<��(����L6�_Ҡu1�� [br�( ��A�@���J�^p���l��'��5��-H�^�+�}����_��kso�.B�d������R��M��8.� �����)d�f��knz�ˉsǈ�r76y�(������y��P`>/I����I&աx�{J lV׮�:���c���L挊���rT֘hfG	��h`���97�$2h;Ľ{[@~4�S9�g���Ee�5n"���sx��PY٭�f�ɵ+	(dDq�s���k6��|SSؙ����&�|W3�c�π��5��[^)}�[{�T/����PX�L�lk��/�ʞ%$>�jim�C��15���/Y��'L��k��+'-hLJѫd�D�=�����I�P�rN�Ha|��[��a�F�ګ�J�l��m�2}dBR���a�u��}�)��賱�]!��B�z��c��]2�+�Um��m1�KYU͐n#�ԫ����)���YJ���Kt�3�'9�#vҸ�g��+KkBc���F.���ZLF����Յ�p���?�
j���%�=Bo�]޹��'-�B׀�><�- ���M�C�1@xa��Kcm�{HU�/iWRI�k����)�#Ǳ�:q���hZl���������a	R��+(���)�#��Ճ)k`i�y���$�����ܰ��K 8+h�g�X�0V��:n���C��r�U�}Z%|������d �Kg��"�ͪByB��6{gc��}l�my	��}��N�a�"�M3�^�w4k��/�ł�e+-�-vN��'���Ùg����C-���ɺ��i�ʰ7^^((��jއ��j�
,N���n�b/�x�(AeA���ñ�O�������NI�+� 畹I�c �8Q��_!��k��ǐ�xE�{��=�����TV�tG� �!c��1�x8\��m:w�
*�f3�&mC�4h=4��>���������^��%��p�dE��u�+":=�m�SZ�o�2�-��#M����
;��z\:�~<�4�n�'��A��\�#�ŗ�M�ldE����cƢ�B� � ���wR`��$�`�����˄ڣ�!V/�ir�Fcs>ã�Fl��MI���P��`S��̤A�w<�`O�vB�ps��/� +�H|�H�����%;�1]S]k���ྤC/�ڧY� J�V#��)��
[��o���iJO;�U�S�H�z���L��ȡ�A�J�JF�"
����<���f�6}��Pۙ�ۅ��(�;�����彛8Z�ü�R�K�V����"�G�c�|	\���"go�ݤ��ҝ:`9ʙ�
sgG�k�8� �. ��Rk.Kwyc���������ń�.�/������ȲxXJŒ��uc�Z��<
��Im��ٕ#1�fm�@�թ�}�-Y	��PM,5������A)��Eˌ�4�����%-��b��aX���v�}ˀ�����jܿ�ͧ�$$b�m?Ɔ�M�!��B�|��K2��Wɯ��х;W�g�HD�66��xA��r�d��z���� 4����cE�m�V+�o�d�DJ[��ZmѪf�A�ZFcv�x��!�`��Ȭ^�:k?�Q?mW a: jv�O9�KI �o��x�TeB�u.98��{l��l?�ٜ)�ޠX���&�I�9 �|�dY��K$��L�H׶���k��$?u�����b� �d�N(%�0D��B_0v �v?m����*qh,�+m��j3�{��ج*1i��a��Â�{9�L���V�}XފL�U�/c�����Li�l�,�����I-ov|���1��>����q�NF6W&oBS���ř�K�Ό0C��fE����������!$��yxH��;���(y���mn����7"�Xz�9G�K�`�t�o���`~���r	��R%{D�(1|�S�)!f�)�EԐ����Z��@�5Ǧī�#(BV|w�������vG[��ӫ#?����#�Dnֱ%�^`�܌r�
���p�ʼ�<��A�iNo����{Z$}IO�_�+���ώ��M�&a_��q��2���3SC7�З��7��O6��׭)bە5r�u�%��W�l���艪�PF~�����7Ekc��!�e�����܆�����ʤ@GTfR�8���`���ֱ		6A��h��3$�b36��p�vlW�1{����>��_��4�R�R�_b�Ԗ��������DE�O^7���pF�A�L�;^̬�L����d0?�9 JdTCRູy$cm�Qȷ���S�.#�[��c�5��o.>�2"e�1T��j���wx{	���a��u�De�C?���N�ej�~>��|�T1�<3�B��{��}��\�_�������X� ��SۑH�H('��	���� 2���5`�г�dZ�aح���!%��
8O+.��؅О��>dǦ��B9��bsj�������� ���V��>=X��N�y��yi��H�4=���Ӻ�gr���u��'S(�;4�y��"ӃX�h��=�
�=��ִX����aa�FN=NO�Լ�V��Jѽ�^ʞ�����2�믦��"�`5�b�JC��nW��t7��� �/K�I��^�GN�)��bG]�2Kw,���z	P�x}.�u��;�Ƒ��m�٦�~�G؞ Ϟ�-��*p��+�%�j�PN�zT�ԫ��Ի���	�_�ۮ[O��,bA�1]���`j�؏{{I�<��Ӹ]H7���h͚���J_�{S@0]��C~�d��E��7?)���r�٨�m'_�AX.��d?����ΜYx%��CKG���/��q�b��G'�u>#K?4��������Z��1=�b`�R�Y�}��Y��Ъ߽��^��w@�$>TY5�Q X�Fe�v$��cl0[�&�W�D�u!�r�ɕ���~ @3ʢ���3�ѣ<v��X�D�R���&�7h!��n�Jh 
[/%Z�@��U<�F>��t���N�:& B!;5a�I�^��isܺ��M
Z�ѭCR�Ғ���했�!��Rnj��?����i���f�^���@�������f*�?N��	��/_��h���4�&-�^&R�R�{º��b�T���"�ź@�g��B�b��T�LEXoP���+��ڵF;ٹk�V�w@x�J�$��?=�,����c �����ի�{޺罚���6<E�Ͼq۰ŶZ���B���o!ʁ3�<o�2��Q>ۊ����H2S}	�57d�%+}n�a�$/�C�}$6g�!��騫��!T'.dN��c?#�j�kg���Q���t��tq�Bs��#��2���AkOw� ��٢��}Q���jv��ƃ�u���F����z��g[ũx�CR�5#�F�x�Y�#� ɻN�ӊ]ZHK�#���J��J�ٌ��Vr4��/`=�↡�"�p)���1��PH�<
�ѭ�ǣ3��@J ��L-�@'?l�
O��t��a���%F�Cҗa��q���]��	v�H�{s1�x(UQ�"v�x�[m��/��4��� V
�/%�'����Y�� ��"&V]�٧���˷�d_n�#Q��
��Zy)
�M�Ϯ9Z�K�<� QU��f�4�������I{���PQ�x��a,)�U\
�l�.͠����4��޴�+1���q}�L>l�onm��}�^�����9�<��!�c?m#��
�cZ���A��m�`|3a���u(Yu&��b\^V*�7��!��4��J�C�A����A�9*b**�O���4�GZ�{�K r�i��~y�pEP:~<S�����i+�g�TT;EQ��2Ep*��^M�"w ����E�B
	yn�)DV 03�#
��J�楚=�S����҄���;��Gr��6�����[�.Է͈>l�L�[HT<c���ݩX��X�*�-lC�z&�$��)���T�Xf���&'�_φ�|�!�K��/��.���:�Z�I�{�`a��9�+|_9��Ej�a�}ҿ�v�0����G棾�h��]n˙���L�/2�J���=�C7;�̢���s����A}�8Wtсm��~��k�L�o��b��٢(��(=�w �ʄQ �vȀ��R�6�qG�c�r������t��'8�����T��@|��<�4���m(�����
bv޼8��h����Z
�:�p�K$o��g��
�r�<�s W�8f(�h���!�7;�!߄��K|�>50��ӣ����qZ��K�i�W������J,�-h��TYO\~�L��?l"�7��)���
�_T-k�g�� �T���J�Q�6�b�O��4��0#�9'��"�iAE
H�6T]湋%\�l�������s�FϼvÛ �0����|0���9�=�As`	W�?S�Ȭ���q<|vy�2��Ы~6pf���on*;ɑ�ؿ !�iH<]�YPMh�tw�� `�\�3:��O���-I�79/@q1�1��m�MF�0��� ���Uy���qQX��Db$���j��ђ�	����̅�X�E��Su"A�@�o�A��j{=�棢��k6\ϑQXwM��'w���&�r���F;���P�.�ϖ��)
��8�4�'�~"nR��/�K%G}�:���ۅ�xE{Q5_�P۱�m[�؛3��z��OO��:q���))��|6�ǽ�a-&
g��
�hSq�~y�#�:!il���>��/�=�^���C�S�������H�>7Cx���zRQ6���֟��	ް5�%��N�3�I��@����5�����B>���;��� p�pLCa��l�ȟ;G>e���U�$�v���z#C����Q��lT�"c{�ᤣu��.t�X�0� 0k���w�?�+/�J�*�C��s���Kc�U��84t����{}��j�E^���e�0���h�SPݡ���NA''���R�YN��h��Vƶ�m�JP�r��h��R9F�,���ƚ�J׼1]�.��LY����ʃ�O����Ĭ"���~W���0�h!I�픚����?�m���a;Q�+���L�.l��̯2%�v�ʴ�58��H��
����V7��x�8T��e"����#��Aľ!Y(|/ ��>f=���/̦��#J����l)��}Fĵx)��G��M甑�7{�������!'�F��E�f��x>�rT���/_���'���`�> �>��1�;���H�V�)�d1�fi}����)kH]e�s �6�jh��	=9`�
Q�AoF6��*(}�r(����wG9]��_��P�`��cx{ҁ�cu=4��ߞ~_��A�p�L�24��*���:n'��"N!���PO3���_�G��;���������R�Ω~�Uq��7��&��\,B\EFW0J9�� ptMb��(�7��L[�c�f����K��"�"C*�J�]���x?3�z��zn 3%��k�C;uq��@lo�����I�rh�23��5�`笑�,��>A@%��
W��~�I]�L@�����(�jU��zH@_��ͬ ����o�X����>�k9=dS_E���N�ˋ����� �<ڤ�¿l�)+�b��[��&�����6�l���[ID������0�۞���?<g���0��]�;r�N�q���U�����ϡK�Y�H���_Py#�5׵�\��� (W{n$@�J=�*��u���L ��D����57�bQ���T�F���𓑌U~߼�ߢX5�J��	��p�'����N.�}\ظ-��g�\:�LM�kE��G��6��q���2��2��`�"��f��+yY4�C]ɥ�6�ڛ�F�ӳ�>��6�VӲ���|�����~4S��ͳ�0��*����9�K+���M1o�Z�(Z��Q8��������U'p��Y�2@�=(��M����L�: ��1U;�e�'��t,���GL�z��p���m/z�P��C��ݨ��(}���emЖ��nN�C�3Tw��r
���ކ�I'QjH~�(�x��ݠ��xب���Pf��M�*��qm��O?�O�>q&�;_������h�R�2�6��{���؟�<%L'����q���ѐH/O���=6�K ��i���sY�9Z1��rp�$͆���ǱN�����j�Fl|}����W��lO7��bwT�����˴k4��P}���HB�Z`4��G	�� �ܲt6e�)�U����6 ^
ފ����$Mi+G-����E�����fJ
�5��r�Gʘ�kR���H��\A[����>�\HJ%<<���}:C���f��8�l�0�A$W�$^&�*���#:Ө����.�r����!��oA?S��8Z�a~�g��K�#��0ۡg���.�6��z3��0�&e��K�:d:2ۻ�\1a���sH�L�E$�J1	�{^f�3�2�#�gI����@���/�̱�*(bC�yu0�%r��8r�LNރ�����MQ����V�GHOewJ�1�@�������.n�ZX�~�N)�Su��]߁�we
 ���NJP(app*����9 :�^�Ԭ���e>l�_Zu��8~�n[��V�ը| ��K�"�۾��D��qU�����F4�;'���]�BJ�ӂ��6"V�1�,yI^M��d.�Gi�^�/��	�b��|��>����N��,s�20�����L�����n΄幋A��.LK���Z���K���L�	)���,�S� g6�_�z&1��As�FN	����Д�&�"�'.��=<�n�a�9i)�%u;��!�9��L^���@F��Jۀ��E.�Mg\�{[q��s`�L$�Z7���)���HjBu��'~ ��\hd4�'��V�&�	C��?~��x��������/���Bj��¼�)��d3k����&^�vv���h�*l���33���[Z�By��DEGk��
��-�;����M;��<�ISJ�r���t�f�[�yc�a�Ov������w��جڀw��e�?�!�T�k4��n<Z+gwo^�i{�%�w�W�(�5�Z��޼�?�ԉ�[����>�r���p�P�p<�&80n����(�-K�m��F��9����ñ�Q����؃�O8�&��U449�P�a���L��ν�����԰^��,�1m��\�$ ��DӔ9�=�Cu-�Zf&ErbErD�w9���3Q�D���J=�!@GfO�o7/���`�'I�K�i��`�5���f�4O�\���z��6�h��׹��P��M�c�0CXb:��\8 ��Y�b2����Y�^�>jĿK��w�!'�5�P��A���.BMD�m�v�[��%^X��
+iI�ሖ�,ݤ��k@4{T��՛����W�@�{�Ռ{<�����:͔� 3/X;��p����Z"���6���]�rոL����o۫1�m��p	�n�LI��5!}3EU�����"��kc��-��Z0�yV�w�R([�ڏ�2����|��g#�-t�{.pA�B��)ʷ��  ó��m�ܼ�~m���&�+���1�+GlE�&��4�ɸ�#��ޏ��@pe4���M�A)e��I�~l�M��:�/�ѷ�΀0��k����pE�@mt�Qz�_��,8�x�J�WY˚v9�����EP��+�"6CC������k�X�Hß�C���Z�磔��v�o�N���F���Z��"�;��i@Y�X��S�ѧ��쎪_�ȉ��xի��G��ޭ`P�.��5��h���7Zm`c=s��q�-�(N]M�Up�j����j���p8��0_�d��,ׅ�X ^srZp�Jd�)��ɟ'���y$��q%������#�M5�?r��!�UY��MBI��A����S�D��m�U I�8M�HtKeB�TBL��}Ӎ��Hx%H畳�p1�6KrJ��>��	K_ ���.��t��{jRR��u�5��r�:i�X`�IpY-����O��Ѣ�8���[�9��.�YjH����Hs��E@���3�o�R�@�Io��@�&��Y\���z���yn߰gd!����F��7[dL��~�����T���<��z)��i;�Ѕ�������T���<
���i��Od�L��&��P*ȁ��5��4ݍ9a��V}x�����X�=�G�X�R�"��nq��]���q�n�o����Lp&F�)��L��=)�~�j+����&��Z��ֹ���1B,��꥙�7�[fb�#)�+�O���HQ���&�����v9ޚ�N��uP�b���\_�Ԯ/&��h�u?8���b��eƓ���ޒl��GIt�,�g�g���`,Ie�8'��=���{�<��M>C	���������:Lg�����U��#��J�'T۷��Й�ٝ�V�tr�~��)6���l�oy4�]������7���&SMP�X����P#[�d�!2�
�l�uu���ñ!�����q�� ���<� �=𫂫�^��n는Yw��j!��t(�Ҽ���MΤY�}�t'f���P=+\ 7�l���T��D�]�/��Ƅv�$�b^�x�����W��9>�w�6Մi1%{��o��?K	I�ے��;$w��W+����_A�7�e�d����d9�]76H��@Ԉ��c0$�ܔ�&r��M��V+9,�-b�>)k�1z�l�5��d/���\�P���!����U������L/�KЎ��c�|���&?OU �wGw�>|H��fp@� �� ԧ0�9^�ܡ��=8��v��&�$��&_T��т��q���Au��jHY�\\(�s�?O2��- ��Dx�CMn���W.ɰ�^��Z�k|�=�;g]����#��ͭ��K�cŷ?aآh��+�Ы]4��ç��)b>7L+\ù��3To}:�5��8�c?���PH��ֈ�T��ڞi���Tl��1&B���X{ͬ(�*�B&5Y�ϙ���c�R��P��@�,�j$��f(��
~�]��,�.�T����/ъѶ7+��n��F�5H#���]ሦD�d�Q���vo�@[sJ�����l�H�N���.{�[��j�U���%=�Wk�NT䙲d�_9�=��x�1�/�Z��Ӈ���Y�>�֚ET:�/t(������&�s���{��@���(,��b���>/�*l��,��Jם3�8c�(]��qs��'�+"��8ih���@��hO�]�imx!3`�w���JZ���Z{x���� �MCz���Ւ�)GԖ��$�:�)�+W3�0�n>/��e���EMۯ�gI�fu��=Թ%ҵ��H�7T�A�@�>�n��߈$���[F/j��C8