��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F��J>�����>�����HU�k;�� �[�+?�w)݁)��>7Ý�4�B#�"u�%��R9�*2�	φ�v&�f�UxJ�%�����OOL�mF4O0��%�O6?][��W5Ff�i�]�E҅u#��Vg�n�����g9�#���>rh�W&��zCu�M��{����,l6�`I��3����
X�	�@�#��꘲t�}p�ũ�g���.�pæ�dbB�:�`�(8����Q���E�m5���[\[��Z�Xe���z��e�ّ̀�4��'͐??�r���4U��e|{��s�_
���^��5���ЉS�u^R��r	
 K�Ԓ#tO���?�M�ΟuD�(}�G���|E�,n���;��"�z���+�rW�t�ǟ��[�z���Q��Ƈ�b]e}s�;�H�:��(�=����ݺ�����)%����j�⽾I���G6
�<=h��/�[m�S�\I�.4�A�1��S�S��h$��Mj�1�~�P|ul�P�,hM����R2��U�&tˀ.?���9i|������u��F_8�����-�'zx8�~�$	�	+��D\ߍ�b�+/n�f i��O>U�9���mx�������V�K�`?2_�ĥ�3?@A�ʺ*��P �j�C�
����ï��b�A����[���GE��\
���k:
�@�fv6�xR��G��� +�U�.?�T�:y4�_,��7�&��!J�+9?[X��b�1�#���l��;�l���@�7��-�c�)��(�E��V|��i�P/��0��9���E��bQgb
�fYR�E���Do5�����6�r��"�Ҝ��9�=�N���5�Wؒ4��P�bЊ&x�`
'�97^�(9�!W���Dxp@p-/��0Iﴓ8�Y���v-qk��;�Ң7ժ��ٲ?������TH�A���o~��pI��<C�@}|ل1�ў%hz�&��-p�n5�,I�)3�����*�}{�.�O� qI�naG���"0Bσƥ�pl?[� ���,.χcFP��&�?uP��
����������K�,��hXJ��Q��^�M����ϕ��< ������h+ycmh���I�s3]��6�  9UĿq�����⨼�LKU����,��#(w����[L�ޛ���N`c�c x�j�Z6l�iq�ﴌ�P�	�:M����#Mt	��(4Tq�4p8%�;� �o�;*�;OI����˲n��>Yb��EL||;�Yź�>-VRx^$�S���/�]��{n�BX�'i����f��#��:^�:a�:����1�./���)6sm{z�e�r��?f8�XP�796��ߑ�]x�jg�o�۟�­x$_����L� 㲔?��r��t`j�{Z^\�L!����k����S�{i�z��n�ӡt����&��KigS�a�_w
����Fu����oe�k�XVM*E�pbϛ=��nۼ��"Ep:�����*t��Z��k i~#.��`���A�ȋ;�u�U���'y��ʚa�8n"�f�&��Wqf/��D�4�8nBmFr��@���������
��|�QM��<����k�&�di|g�ᄌ&���S��=1�'�:��[��u�b7��jQ��ݼ�@���E��k1R|*�뚩�޶�(s�.^Z�B���"'�dk����]*���������H����H��M���LL<�[����e�
"(�h$)&�����Yz�-������Wb/�H/��<�'�Z�L���2����q�LL|�ǖ��0�q� f��!86G�l���#S��G��˳���[i�׉� =��E�]�Բ�}^�i��z_�ؤ�"���������;s�=�o�W��((�h�q%���T���-l���5
V�$���e���@�D�N�2w�Kх]�6ʌ�(� (�W{Q�x�Mf�EpeÜ_�)_3>qM��aR�ɡR�:�HDK,�#�hu��5�~�����⺰�Zz����:��Fӥ���mL�&� h^�͞�M93�mh|��C��M��o%��.FɺH���p�Lz�/����[�]���X����Ae1�/_���U�K*U7?�6� `�Y�ԟ*�k�OJ�����3L���ĺA#���P�B ���C+
䲑��;iN���A�%s�<ḙ���=2�h�o	��R@����r싕��[\A��'cq+��k�� ?���7�#շ L<5KL*�yA� �~i�\���D��Z�ǜY+�j=�%P ���gy��
GR�HU���I��gY.�Ǒ�Cs=�HW!hV]�\�J}��}O{����\2���E7t��ϟ�q�\��=L��hQc�v�
��H�U<�����/+���S���v�e�c-7���Cji�-^��%7E���7�W���N�pA���I��}���p���dY]�Ƈ�g��d����g<�
C�Ǻ��ͮ�.���;�~hK�}վˊK�A�^�ah�u��"	�O��Վ?� �5ɠlR � �lgo<� A�_U)ƕz��E3b����bn���.W��QhWK�A#�:�U>��g�
�DR��]��`�|��J���#K�� �cj���O��L��|8�����q�U-Z�#PZk�5ײ�:k���tP��x)|�®���6 �!t@m�Ao��<�A�.�s&��!e��\��x�8��i�6n�����(�Ο���V����/ֻ$�`�Ҕ���� $G&��aKD��-IHj��� }�L+�0����oi�W��vLi�͗L>L���ɸdol�q��A8j�+�Pآ����fC1N�	��/�=Vn�{�P�58쀲���$8�W�:Yl#�kX���ڿɊB_�ڮF�Uͻ�$T����z�@9���'<a	��i���)H%1D� )�6��8�Lu2u
�{�[�k���
ߘW��irM�BR!?�p#�	��Sx9��53;����h��i�饧Y������~�zA[�J`��O�:7m�Q�°\�����Bo��Ohi�d�(�A/��kw.L)�+p�K�u�Ƙ��@H�1�����N�m2�P��x�t\�.�&�puĚP�͌��R!��5�?����!4I��2��&%1���{��e��C�ԝΈ?��o�l���Xٔ�ڋ���:7#�ڸ�" W��'c�ӄ�h��'_�.z�Ϙ�1�d���T����+�q%�?�Zp�]t8������x0��N�M	:��3/�wz���L�&D��?��D01���ϙvIW�)_�F��F{���Ҥ<G���T�P������Y\�)��s�i�{=I#+M&Y���!"}Y;�J��z�܉��e���2�o^i�X2���_+7.	�^����P��3�t�r6��]|�ד���xC��0�o�̎mи��Xf��d�y�'�8񰤫��<�V)U��9@<fv�4V�QE�l�mT��=��E���UG��r�1�b� 9Z��e>����F#$�z�߰⏝^��O#��IS��cք]\ĝNH�d4۪�잼��B�Z��L6���x�M=�5�������������E��=daq�q��$x�҂�d�@��%<����	�y�vD���yqCdvu�I�>
V��6���|�m��הd詉�f���ԥe~�O��-���O �����$�L������kC�O��edy�tH���%�N�놮'z�Y�,���ᛲ�� �
�������C�^E�_�b��BK�ל�{&�Gt��KD���и���m����Ny��U��4J�l�E`p��{�'�Om��d�<��=�+�����Z��`�\&V�ͦs`ш獍UR�[��������Fv�֓��K�h�V
jK7�(D���l�.	@��p�9F/��b����uo�,V�L��\=ƛQ� �ԗ5���G.㱮�p�߇��l��jSe|����{�]Fn΍�m����|�����E���zR�')Z|��S)Y5eD$p��M$����&�.����p �[Jܠc�j�u��'~]	t���"���Ł��Fp+^�5:�b��d��:�A]D�7��C^��~mo��_|�\�̔�'�+w�թ�I������^M�J&�����/vQ*2YS��4Apk&���@�)��c׸�"]���r��q��v�o6��*�I��W?����EW�}����Q�yr�~�,�竣+�.�E'�vjC6b�x@�q��{��g�r��Mzl/��
�B�`cC����Ya�w���z7��!{�G�X���Z	�]�}bQ䔺jk�3,
���?���A�㲈.����fDC)�k�����tݠ� <��0���+g���=�
<�U��CA�m&�G[Ck���،�y�������3�#�D��<��X(YI�b:���0��A���13�Gb�ك�2-�Ng1��	���,ܥ/v-K%�"Z��6���f���հԋG-5m�g�؉�Ҭ�ڐ �td�!5�E(.᜕0h,�L$s��]iH6`�8����~�2z�^6�����Q�zXuu(|l�6zͼ�0�:'�낾��W9��\�q���g���O٠�n���|v}�商J�X�������r�,�]x4��b����J ,���B�o(B*\�/�iD΀%�]�8��_ӓ�I�k�f�!��5 �>-��������]���F�,	�1-U`��T��ۉVR��#��<e�'�g�	�8���;�~y��Ķ�iа��>��ԍ �5�p�s������T�����\O���o�[_�w�ǮȻ��q��U����(#��GP��l��`�r�#I�#?|��g"]V�"�0/$�"�K�Y.^������������[�;*YaA���޵g�Y���0�!�X��h�b���t_ѣ �>DIMz����\eM��@��]�^;��U��L�}y��[���s.���a8^��u6�'۩�ȏ���^'qz!"ݥ�G��R������"n����ZV�R�瀶���Z�z׷��0�������������Xl�wi��~VK�[#v=!�2ps����A�ʆ�=J��f7�6尺��vυ��̺�^��s:���͝p�]���E���KQqL���'ӓn���4xR������Ź�$�k^MJ�������F}TbFHX��>�|Zr��z�Xa5����z敺�Q�[��T�?&G�ltЏ�bpɺS�<p$ƭ\�g!�����鴒���5��v��
��]߲�ք�/�P$tֲP��p2 ŉ@�,� ��8�v�Am�.�%��m^k�F��́Nb�t��?�vJ�T*�̕.J5��w"��|�AËl���\��:6�kp��d�/a7߀쁰	���2��씲��QQ�#y�`1)l��!�!���x������Ȼ�kQ=�h�"*+J�d�^-�|�+!�^LL`x$�Z��4L���֊y��h���Tg�Q���οD�}M ����c+߬-`�$����J���|�i+���1�7rTG�H�C�P�!�����G<��������	��\�j������g��Ln��)Uy;�"}��1���^8���npY��2�>�Bc�����}�mt�@��.��J<럧/�5��Q����4(�֟�N4���|&��6���s=�:5���'�b�����
"dJd�K�yQ�~���bWL��s��#��4g^_[���"�H�Z8��%c�n�Du�ы̽����iq���b ^�iBqǡ��8�ӻ*�NV/Kz[�r0��?wQ�p��<�1��9S1l���j>�M�*�H�`����<��n�p�Q�I��2���	�0���8�����Dm2��,X�χ�۶Dk�2��4�)��n�|�^[��������n��u���� ���f<�8F9��rv8�:���~0�
K���C������$�\���E]���-$Ea1��&5���L�op����ʮ�����$���Ӽ�"ܾ
��.���N����X.��K�ꟌI��ޘo��K��]��x!�4͔P�;��;�c%���!�t��8����N�)��iFV�~�Hn����Ǖ�Gi&�{K5��W:!>Y�4�D���v�_�Hz�r،�f���K#Vz'OG}xm������T]I>�8S*{4�t��Ps�h]�c�ݹ����@K}P-N��A"JW������Z�pj�n�Ŕ�u�bc�IT��.X�o�c+��5;�_�h�}��.Y�y�.U�S�i��/?���Z�+���륃��C��Y@"��grE^����mI�d�O�F���oHO����3eIuh��
��w�=h�� �ƢK��,�g�
'.�JC��3(�!��̎�;�s�WZO���R08�� �o��cl79ܘ�U_����@k�E��*X��e�Ā�
ɖ�l<��i��e����äup���{�3Ec�v�J��{�X�?�!!Zŗ�d1A�R��N��lj���o�l|�
,jЁ�.lP��6����!��
�J$��"��1��^lR1��QP�g��Yw{��鍖O�����U�J�����S_RC]�"�X��s�C�9cIW���m�i�9���Gko��:f�1�dSƏ=61�1w_T�×�J����aD�H�$�BP�����w�z*�Jy��0�s�,}��o��K�3��D����<=.4��`�Ʋ���hI4��)y}7���5~���(��ם�����,�|�ȵ�#[�#NG	�,����G=�M��2��=�K0��T�UHD��Fڍ�����V��v9Y7�\c�"�4��q�"�i����ۋ�Y�9��۩{�J��P�s�94�*j��5��u�|�PUpB�m�P� +n)V&��%�ӷ�����2�`��t��c៤�+�&��v(o�G�Op$�����
r¤�o��}���d��k�7��ӿ��vT�,.�xE�0��C�8�$J��d/g�t[ �SG� ��d�!�I����W���a0��K
�T7�X�x��[&�4�$:��,ʑx@����Q�͕=lQz{���|;�B�Y����GK���#k[¡�"�*����z����;fz��H�sOXG���4�
�����l�m�A�".8Yq�BqD���� C��q��"$]Ɂ����dݷH3|&+X^��:K0d��&GG��D}�:r����%`b���z��0rgvr��܉�/R'w7��$X-�u�V�yy�J��bm~�R�'q�����.�'0�^�ԕ�Q����g�u��K\'����1�g��K�����]�=�̎H�d��k��d�����DJ0��u����hE�X�爕i�%$�8`U/��[E����f��G��~��*c�����m�7(��`����X�i�j�������N��UJ8��q&B����
#L�� q�H}{�UK|��\ |Ό���oH�,0��|�p����NQU�� �IҼ��뽇G���U�v�-��,g6Y1����W��ڃ:�"Ǻf9��%�wT�X�'���˂"H�\����H�NV;!i���u�)z0���a�ia,���N��������|�.>Գj�WjB�m]V��a<ZU���	�NQJ�����E�Ѫ����O���������/�o�}���={�A�I�ܰ��h&�c����'�wHt�p�mC��:|�Q:w38+��q;�r� Sg���1�RC�F��?f���4�d\�B��t��*{0M뷰L�n����V�$��tv9� �(<����.}�r��)X�]y^�3�a��e�@� )�k�>�#ـ���J^�X9��v�d�΄�.�ֿY���c�c�|��f/���%.2W>�D�R�[T��_����'W5�d��T�o�kC�B�_�,����N)O�T�4��'��1bz�Bd ��}~��u�i�H�r��z�I�7�p�!�JE�~�^>����&ۯ���c�{��-`F�#�x�)z����#��J���WH*[�s�"������u�vͱ�ko�P�)����FA0mŢ�6t�0���r���Gn{��$�s��@�Ta��q;�W��=��[$�ָ��@����nA�ht��!"�3m�xD�P�RՅ�9�la1%̯�(4�C�l�|h��ih�?G��(v��[��k~���=���c�. �kG�\Y�R��"�O�����g,���Cm0Yk����=����H��g5������xk�O��O�L�d����
m��]b]qi�=��U�Z>�M�����;��p���kQ�������6�-�n��	SˊۑH���=k�"OO��8X���Z]�a�k��J��2�	Ha�3?2�7/e#rk:s͠�Uq6t�1Ů�;�������꯽:00�XqAT�b�O?*�._�(�5�C�t���̜٧���r{tѤ�=`�ZVsk)n!kkk��񯩕�;��$��z��@d�pȔMVޠ�a��#���u��IC�mSS	�U���ǒM�X[Rؾ�~�����;6��8C�9�=bh��᪉�/�1��c�k��H�+��2r�w�i�4`>�FO~10Q^(�.�l�%2=�~g�i.��ߢ5�^I
E`,���	��l+���|��)����O�X��^S\�d%��%p
��0)���r���Ϻ?7�e�ő�i�s2���!칩�އ�v-x^��$G>?�>�-cAn�|�AhQo�elC�W,cC=NH��,Yg]������r����k�+�N��JbR��)� �߂U.���l��i!�C�vS�.�Q=����v3J�ȃ{&��7{�@b�����~x{'QiE�&��������t������*Qo����v2&a�E4�(��_�DM��[��ł�s�p���0\�<
�\y��K���}�<HH|V`����yg�<����e{�Kt�gV����g�k����ĵn��"p��͞藃�1(qc�51&z�e�eG9�k�Ϙ�½G�Mn��5|������O�\��tÿA�b�@�&���I�TY�$�Z��\�h�� ^��]qrH�����ȳ9-ȇgldM1eS(�!`�q�Re؊=���u�k�g�Z���>`�:ȿ�����č�p�U�@�_���+%*o� �Ͷ8�p�hBwh�X�z��P�M`Uri�ur��}j��jkx+n�돘��V;�(��r?,L��t��^ݰp���5�i#����q��8 ܡ 9�o@�d��:H�'W��d��`p�2ڕ�-����?��V?�z���R�Q�ٔ��1a}kS��u�w���i������������p,��yo�+�''� G��U
$4EPU7f��ʪ��.�Sp�a��	���`%����d>�iU����^H�}���V�Ռ�Jco1đ�8����4��|�$ߔ���	��|��v�Ճ�76Q�OҀ���ʓP2N$YE�wj�G�M��Dߙ%:4��<骋=$]o�?��k�x�SKۏ���څyQ���2�D����3h�,Zb�(�oO���!��C\�*���4��a� f��)���T}�Jg�*Ŗ��N�5�Ӭ��=�z0����=pbU�:,L���(�s�v	�hS���U�ȡ��ҹa�o�(�a�&-zhk�s(h����<sԘC(]�M	{�(�����zF:���&[{��4<H&�I�Cʿ<���C��_VN.ov@���plc�r[~��:����:oƮA4J�%�*?!�����#�&�D��T��9���uj��3\���IS/A��E���[��lSV�P)�K
Wp���Y��3FN�8&`�ק�� 4`�r�7i&L7?�Pˆ2�oȺ|�1�r':������cv�١��@ �m9&Y�C[�|�%L�	\�(�����N��G�pVnY��	����>��.�D���\t~�L,��n��;*����<?�{q����N]�?@}?N�3���x_����|��S<̝j]�s(g��|qE8��Z�4U�#���s#E�W�bo✒@落��Ĕ�j����ۡ7yU>Q�%��<LT�+z��c�ϳ��Z�E�r����P���z\�:e��0����	x�T��oɜ$�5P�i�W�k����e���q&��(.���l�8�ﯪ�khq���H" ���o��q�N��)x(.���xh�[+��Jf�A'u����`�__�z�/����ˎ4G�r�C}�|����Nt��`'b�����G�85R���v�m�� tJ)�]\Q��
`��"��y���r���h�]�w��՘�������C�3�L�w�W��d�4��_���om��n2Rr*hV�|cį�E.=�R{�{>lm�����ƾ��y43�A����
�l���+Re3�N?9�7��a�O���᫪^f
�^p������V���]�ߌ)x���@�w���d �����(����t��uGSo�P��Ά0�dO�I�;K���Y��z��]���ljB�g��A���I�(ٍ�,y��� MÌ�'�^��U�d��E�`�I��7���d�P��	B�|��f}�=Q����ɞ3���2�Ĉ	\�gy�J�;���gz�k�i+Ӯ�����u�l<U��Ҙ�Mx�*��~շU}�mJ٩Z���=<]�~�/���_j�jW�7�v�����I��Se����Am�](C	0 �ik��'eA�_���{�p���?o��\��0���#���������j�=�Ė������=�""M��Ҋ��E�j�Z��� ��$0�D�Gk�(ʘ��j�rЙu<�O���ɘ}	a}E�]�B�׼���pS.�_����
 RVΆ�u�?�oڿ`J`P��e&��6��W'�՞��4��
+���z/�!ꎵ{I���̚��s�M��m��pϹG>�u���P��>d!��-I���$#& 례�_K�fm!8a��U��_�����Ǩ��L���&���>�
s�������6°t)��r��m��4�I�#�;:�c:t={�P^��7`����C���=��a6^���x��(@Ei��#�=�b�Ee@)Ax�樬E-�� �8���t��!�+ޕ�޾Q�vAF��;2��d�Mq������9�68
�^��H|��x�4�ps���3Y%:��X��52�?� ^+r�����i�;�v��/iA�]�3�ˌ�8 �"�11Kp����c������n���U�"*�<�k /;w�z���x�z������7��X� �y���%��괹ޔ��4�/#�	��
�����^ �"<:���Zu!^Ѹ'y�c�P�Ү�j���es��ţ5�����^��`���eQ�5B=�7��Lhx�T��ﮗ�~O�  ��f�<����5�+�� ��o..�du��">X/����x�A�r`�9������]m��F�?S��1��l�L�UYo����^�u{4�+Ȭ�U?T!B�+L����� ������s5,]�Ԝ�^J�08�m!��*쁸CEۜ��+*ƪ�M��(��b�X�b���u�)�͵^-�x8�9�x�����������d9�}(Y"���E&�ʐ�p� Y��s�G�oQ��*M×af
�"�zPt:�J��n�����ymYc;�|������x�1�"ۅN{T[w$����_�9�;�1��:Aи��;�S?����t�kO(p:@�����U<Hi[�g���"1G짘�)U�
*�]*�/;�ڢ��3�2����rR|:T��k��|���s,^�R�䣰y�g^k�BAj֯l�)�5��~����͖6<<I\���in�/���\��sG�*��C�׎Ӫ�&2n9ɮ��J����޺dv��x�h��{�@��GB��{>�k��Y3���x�p]
W��+�7�~H�a<S�s�+��>��K���	,k%V$��l"{��+@-|�q.V"1Rv��E��h|��y;�7{*��ؔ<�Txp���wL���A����Dx��l���=�@�)��HI,�.��Ъ�� D��p!�(C���s�f2'��̂4��!�� eF��ؙ�7Xb�W�SW��ڎ8c�B�� ,�����7�S����;�T��+rNsȟ<�[�#��Gю�<v��S:i�11.����7@�Q���n�&-z�S��r+�B=����]�3.�q�F[�h�-�L�̎�U����u��Rڄ�ޔ���t���ɄʵK��4n��/�����.n�8�ݝc�E�-"�_x�)�f�GԒ�
�xZ5�eB/����I�*or��t����ZԠ$~ �(r=̂H%��x�Ppz˱y���`����7�œ����n�5��� W�`���k�'��u���:�KB+U+��o�ydÀ-51�.�{k��{��q#��
��R�����G�Y]�X(y�.ֱ�>2��?��l���������ך/��,�iZ��OU)���RF��V(��C�A�n���b���&w��)�
!���B��*4u�Jjg�� ���L������v�#�b���_1��0�2�!�9.1lX����5bҦx@�%n�#���볣Ԅ}��=ϰ7��# �Q�	13��^�Dy���[�湠�o�7�`o�C�c���Đ�1��Z�g
��<�U��%��
�8oC��P$C ̎�A����V}�;��3�ؔg��B<��8d��ih����74���!���LX ���b�r�-���� �D��P�3Z��hT7�
�x�<��w�7JiV0��k��	�w�4����+�T��b^�zBy���$�	�z�xdPʸ:J�y����-�<n�,�֊mq���N� X�R������u��x{O��ӎ>x����$����m}��2C�^K�����]0��a��H�2]h鏈t�jm�O%����U^7teG�y/s�F��o�5�n�ӒŲ�9���J��w����g ��f��+��Qp�zwbb��3|�C�p{���w�-�V���$Ƀ����·d���5�ngN��Qvf�%1p�8a�Gk�b������{��o~R-�h�8Q���]7��=�ܓ�o�芚7�t��A�����/�?Ñ%[ڄH�������1M��ٟ�k�+���o8����Yrs5�d%�D4m�(�K����?S�
�("Ő�Na<w��|���QUoX~wS���p^Jo�ϫ�K����R0���9T���N���82�e$g��򠙻X��xЩ$���"��B}c���������T)׀2 �X"ȥ��ݡ���=q����ݔ`�����ONC����y������j�{���Iu����ɷ2�ڹ�&��ƴ��`9N�Q�,\���nةA*���N���	����0dۜJ�-&c�~YFL��C&i7��}�/\6s>[�ACKWy�ɷ�dy�qT���n�K���/����4��M��6BH���'>�h��6x�-��p�۲ɮ0Kuf�2:��s��B��b��>�u~0�,��U�t�_!r���I�������IƦ�O�-_A"�|�TD7���c�]P�<�A4���@�k����	'��>�Q�>�~��m��[F��7�]�ŗ����ŢBs�}��,�ӻ�	��l��"c3;t%��CRl�=�P>�pd��ZpMl�y^��Z$��>hcR2�@E�8�	��1E�%*�� szט������dr/�+ף��1��Ǘ���_������A+��Qb����-���H���TB<���ھ�
w��cv(/�Vյ@jva��_��n��ĩ�0J��w[i y9��P���ܘ�Ÿũt&�$Y��cSE[B'*;6Ƅ��'ֿ�޵���;uu�D�v0�}k�f�f.�jpP�V�,7M�n?�4�$����'N�#�5����DF��� ��kK:5́v2豯`9��l1gux� �X�������U@װ�+9����3|�;�q����7���Z0��0�|�8�(��&��=W΀�R��=�S��BG��2�� 7$�e��H�?;�(7�Ӧ�e��a,�ޛ��}~ۆaOY��*#��&'��=�D;�C��9):ǬZ\�n����E�k��6�f�.\��.7�ͳ2���Zn�`M$j3���S֮��lx�|	C�9
V2�W�`�K]�:9>z����H��m8-R��;!C��B2 ݚr3n��wd�A?_�0$�����TPg�Ď�n}ߩ}n	 �z�k������q��5:�O���Qc@MfҢ��J|*`n��*,s�5f��q^���@�������ͣ=Y��roi���!]��܂7G��!�y/d��(���SD)E��F+�'v��-�e� &Hx�Q�v.���;;VJ��Xm�:[|O/�.(�����!�xC�\/���3W�<���I*�䥆�h�fk���������/l�Y/��W���G87K&,��򫅺����n|�υ��]������L��u�R��U��rf�o�l��%�7��˷~o�?�c�����Xh�"�F�M�]�^��7�J��E��"�"rc�����)��D+WB���IlP� @d7��(=��ID�����ś��9 ��iEǂ(VI@��z�}��J}Ҙ*���b�n)�tn�Z�2GY���Sf��9�D�E@#4O��� 	��Q���V|�@�ҙY����<��^����zn�x<^��w�ұi2mK��e�(���j��~�������ŴÆZ������K6���X7j%�y/���S+#��sxe�!뚝�l!2�)<�-�~����� ��-����fߋ@D�Dأ_��i�[v:6E�(�;�%��[]ʗ?졧	���%L[hM1j�!�i:���㼊�	q�O���O��bL�LD�e��R
�mG-&���꧜i������r(�'p����<7E^>I�wЇlLɐ��Z�z���D����=6��`
M��^z�C3~�[߾�W!�f 
S�I��{~�s׼ �2������[fT%���ܓ�myQYA<�ѕ^.���xQR��s%���`ъ_s(=��B����&~�a'�"Q�{x����TkYw���Ce�&;>����!f�˥
[�`������SI%�r[�*vc}��jG8b-��[�.j�p�9�.w���M(�c�W�֞J��~�h��r�|$���7a�	��&e��|�[�W�٥������D�~���p*���`�KQ���:�l���y���hИNhw5K��:Y��Ɗ��L�*N����g�����C��U	MGc�+Y>�ej�)h��!��(b���9���j�l~ʡ]���T��1r���q��v6�E#�o�i�< 堣0��H�������d�q~5&h��A-`��^T|_��/�U%�L�7B��c�&�Ro0ₙP���V��=EY4�vH��������Y�t�3)�[��wER{�	��;t��%����HLk�m ��]o��Ýꘜ ��nL�R�A&90 �����1��V�T'N11@;3W,�lNլC�R����s��8d�#9G��t����@�j�� ⭖P�?/�V����n�R�����b�H�-'u��.�IB�b�n"]Y<�j_oh�����' g����)�� v�iKR£:~�I�)GU�;+�B�Ҡ��Ccc������WoB��.A�P�tx�� pV<yb���ԝ!��cygܥ��-��?�Q�p���Į��%8z*�U���c7��$ŏ�Z�0��/�B��4!; �"w�΁�|���2���{h� �kf�K� ��W<̾�i?��QlG"~Tc��uX�$O�f���#bm";>��lX��Ud�OY�,-�/k���*�2	9����!���[	�WT.i��F��c�
��K�c�d^�-~���y������uP��\��P�\|�bu��yәϲ�����I6��B��P:�~ Ǒ�h|g���%i�S���iL̗�+��_�ڦ���b��"w��n$�R뼕O;��zۣ��SD��S�I�<2t�} mRe��]�|?�nJ�ᗈ��"5��~LD���	C|aO�7�>q6G<��	��a�2M��
ح%��Pi� k�*"��3���q�=���WҤ�:��G䔅�y�H)�z�f�gPII��v�`�k�Prr�T��2��������>$�s�Cf&�2�g�ۛ�d�TN��1���hr1PR5k��y�kkm3����y�.�=�Bj���jI[��H�Z�O^
��0�
�j��G��c~ܘH�	��>,|� �n��.�����DW�S��2�0F��&���<.
���ϼ�2���/۵��i!���#������aZy@��ķ����ғcTC�o�s4�ʙhN����X�O�b9�z��m�����5���k5}Tn3Vamh��N78�9��͂uW�p8�����K�=���\���YM~ݬ�,m��_�0�aĞ��b"��$��fYH�>nM��6��x���h��( ��s��ޑ��ݩ*XKmY��A��j'(L+*QU��h������(U��`B��N	��n�%p��V�K��G�����bY�`�t Lhp�D��le��X§Մ��+���OJ�I�Z8�[��W�
dL�Lu�ƖH�k_C��r�#�$f�&������2�H:攻��Z������>'�Zꩊ��^�obb�T��	��m篊qw2�C '~:� �ŵ���w���ٌy a�^��0�>.<�y=b��<r�hR~3�a��e�
��� �9f���ؘA��l�#���L�t�2���_6��L�nRF~�I��T�7��l�<m�)�<�е�t[�:�ПoZ�7?�DVXBMF�$g? h��O*��Vd+��*>�q($�;2���+�Q/G���8>�S0���.����^�V�!���Xc�x )��p@�HA�A�feH���� ����﹡�D|��k�Uk�A��5~?�OF����B��%�tZ�%�/SD�����D��|�o�>۩�O�ܱ�x�k�%�33��^I��뙺6��x�f�ΩGBFe�e���t�i \IQ�����x� ����iӋE����ӊj����u2��3���Yi�����qa;"��lh��0�M-�@xi���쥭�&ѫ��=�U��.h��3jY�� ���ؖ��ȟ>�·��I[�6�n��F)�>��2s�~��1�Jav~��S�E��C�7\�Ϙ&��t�a��?n�ޥ�]���57AVI����}�&�Ķ�C#d���e����|�p��H���Z�ֵdI��!b�`�����_$#M� �U�GG��Z��#����]�H�M�NIb�Y
}%e�U�D�h}%.��4E=�5�!��JNi��B�>�#\9�G������>�J��5�/3�U�ǒ@��#�U����/'�N9�.C�Gj.�6��|R��Sa�
$Iޔ
ݏ�"&m	[)���
�x�
�VH$�t��O���D�ٞ�T�Y^g`CI�0u:�UE`�`��	�=}�
M������R�t�-��v��@�;Ne`x#dͲ�,"��܀څ����?�:'�����)�zo{��3C���G�8G>�H?��(�/�,��P	�^N�nA?޻�H2qw������ܴ�޺=�!��E#R��G�Z����\߲u���~��~"�ʺ&(s��h����N��$���d�2��DR�4&ٲVc���0\m��x7��'��7��J�
��v�(^)�^��q!�6�ݩ�/���Q@>4ZF�� M��@S �q1�K�����A^�k+����Ej�m�5����0f?��5tJ�X(�<͜1��(]�<�y#9~騤���������8�:P����_#�ϭ���b��[�"�{�W�p<�]'X-e��;��B�����#��4%�v��Y��dވ}/0KE��]��x� ��n�2���0���o��2�z���a��G�:��>�X,��u+�l�R�2�����r�.�F��qv���4��Vݢ���Q�|{��p��Z�h�P���Lq��@T�?���o���V[��H����%��Y��������F7k��2�5m8��\�z�ɂCWI�a�D��y�(��c����K����d�i�M�D�g**����W\��.�}^׼��D�U,�1tԼ٢z���O����lk���T3����N!q�1�����6�-��`�2�j-��u�g4q���	.!I5I����LF��/�$a�\�W�Mn���~�:(��3���Da��]���X��������X2T��#D��sTB��]f
\c��_�~뮚Bn�ݾ��Q��#��Q�7F��X���B���N�C|[!kR�����J���[W^e��*2L���N��M��?���R�̨psv�-j���E����ﶁ��X��P��[H|��Y-�1�i��B>9'���Ƌ���Z��{�~�SՊt����,�O��Ճ� ���P� vJb��l��Hr H�a�Ӥ%C8�G��&����Or!(u����tN ���)��H�{�^4������*�U !S�-y� 6�=3|K�T���AQ8J^Xh�6����F2�S�m��>G�Ƈ�9��ܽ�C�j��k8�Q�U��Q� ��)�O�ˈA��d�I���S"Mm�2ׄ�;A:c�[(\'Z��j�+z �v�_��GϹW/�� ���_�\�R�$��$=�r�����Ed���pP�{�A����	�'z������+�Js��a��3��MBw��i)��n[����C�A�z�D,�Q�0"n�y�S�e_=�}Lt�'A-�m뺶$f5/0W,1A�~����^�;Дշl�&������ܩ7R:;�t�C&6��Oe�c�����߀Q��6Oʶ�L�kI���$��Y�:�F�նl��������$�1�Y'�`�覺�m��.��f�"p��hc̠��ꎧ`Ц�J�c��&XJl̺��J���f�����0ƿ���NN}�rì��ݱ2�?�u6��
�P��b����/P)e��?�NZ��y�b� ���qq�%�rR=�����Y`�Y��p�&��7Зt�_Rh|���mPC�j��*��	��&���|��|O�1R������/�a��������ƹc��Dx1������>����y��X�<�9%��}�ۉ/om5d?*j�y/D(T�_���ULx����my�[�\��)x'a���A�1���x�>�wXC�j�y0P����T�MѵJ���D�Y��=�׷�F�֣Ԍh�^�1g^(��'�6��XˀC�_Z]�'1?;��`f�����
,�x��S0y��l���h��Z���O�Bf�ߕ��]9��%VA�L�cQQ��@��}��犠q},���ڕ y���cv"�g�e9L̸k���٠ź3�YE�dե����=mم�}����;���ل��:Ȩf���XZS�*ā�����Z��<k���w��t�0�!�� ���j�^�>〨����GA%�{��x��+��+����R4��J���[����xo���3� ���VN�"�c�f�b���������ˈȼȽ�So9 ���M�Ө���Qy�IJ���7���q�Oe[أ|�BQ����y���)ktq��t.��w ʫ������	֞�9n��.��~�)Q_b�LZ�AS<I�37�o�A���۠�]��J�9��;>ʙ�V%C���V�m ��/�"�"׿'!���������1�@b7?�������4��
�_���J$�i0S�gI��J�t�xf�i8Aμ�!!�_�%l�F�lΝ¥��/�*�sw�	[��=�����"�@�ZX�	���ޟ*2�ZU��=|Y����m���.�9^�����L��Hx��bG��ߧ��хn�<Lfg��Qv���	L
 Ʈ�u���[����H�1�Ӏ��zΜ��1
�:a��/l�<�D����������u��yU���K�ڍ+&q��?�ՑP�G�̹�(o~�u���%`��=��Ub�fm�|�X$W�x�^L�%�U��En?Mo���38��=�Y�K��}{%����C�dP��;UdKEҜ�	��UȺ%j�_���sXs���y�~�;��P��SsnJ{eX,��G֋\b �������ǭ-���i�+��~��0GL_��WSlZ�4�/͸yw�.�vº��.�ߢ��K�`'R�mb�� �8���I�����8�P��< �����՘v��u�\�JPB���1���rP�۳�Ι��728��>�Pu����	��=����V����H�A{>cQ;@#La8I1�T�����I�P
��_e�r'�{n�"��{	��~��}:��מ&m������m7���եc�k�����5��媘� �%������u�c���	�APý٧� k֧�҇�%_O3K��ˡE�@@�*��|��a�g�n�Q��q��%U��JӴ]���xi�l��E"A��_��s\[���q���a1�F�X�!���t�Ny��ʥ>mFj�6:�U����b�KF�x�(�_qz�����rS�!Mp�5�U�R�S��Ļ�����ft&?f7af�	Ѯo.6��3jٱ��w����Q�_�;�=,��	�Uׅ�,a�Dt���z��۵-�ƓPh"k��:4����u|�1�X�!��&s�K:����mQ�>����r������#�fل~��C����C_�y�$G+�I�0��H~�CQ�g.��D!���	��,g�44*��0w��Y)M�m��ZOb�yt�fz�o[6R�(��=����y��S0)�c��`F֗3�V6]�!1<�C˨��9���4�W|�q���̅�ޏҝn����#�t���[d�'"����U	 ��PZ_a�1�,�DULA�ި���6�)t�B$܏��	�~��(��%�alo����a��1(b3�>1>�[_{���7�a��(������ح]�����~��4�!���je��@.D��nWVW����p�4 ����+aV����s��׳PE8�ز>��wD���A5����g~o�3���)���p:!^���y������!X:P�E���]�c6?Q��z�Jx̆�Z3[�Q�pA��.��g��� VYq�Dd�\ ���:/�=���1SkZ
��N'"ݶ���$c�b�%�"��#X���f��r�LF����M��i�m��v�!�O�^國|;�+�ʤA�S;,�Ќ+|��G�7�74��/��ԕ��\]8�l��=�p	��;A��_���pǞ��T�� EO���
�(bMN ��В���9�4<�������=��Vj���s�ɵ�x���a������Qo"��!�_~V���̥a!�ne}��z����E�8�<��^����w]J[!��v%��|W�z�%���)7�;!��Ԑ��X���=��EQ��a�(ƾ�������m���`X���nf U�;��Y�ү(�f�:#��w(%�${oFj�~�9"���D\K�n�a�j 	~�a��߽yi{��]�\��]��0�h��^��6pB54�۵�BZ�A�)V�&6�U5��I��5��Iݻ����0'n��wk�����,$�
ҏ60����
�@|�x�$+ ߐB��1崊�,�*9����yj^d���;�N�g��K���g���_}Yc��2k_ˬw�́���d =����l�z�f�r�<�q�7���9w��$y2��<T�䶛��H=A�c �K�J&���`u1�{r�����Fl��(�H��h/W�����v�n�%�
��"�x���͢�����`�Bt?-��1"����^�����K�ϛ�$��^h�:@w��6��89
�ꉠ��֞���dz@�ɰD4�7G����x!V����������%��m��!X�x�5��I��w��֏,m�L��X�����ϛ�+ ���Ѵ�8;{�5�'?�>r$w���c�o3�^[58q�I4e{�@��vqe�6�) �-I��/l���Li܃�S��ᖀ���"F�gΜ}�q�X ��(I��]e'\�nI �Q��.����NH+�H���FEK�S�q�� ��vW�K�gAԀ���C0�EQ�*2i�ԷS�W���ޣ����9X����f�s�]πu�^��BR$S��T�=ҫ
/�drs���lt2����&��s��`��5�ԇI�����%c����w�W�l$�I�a�����Y�LU��k3 m<mn�Mt���kY�5o9<a�.��a"���B�f�T����л��xP�NQ���g��HD[y@��At�AYz���&2�w����ᣏ��[����'��R�9u��5��dX���Չ�1���F���U�{��瘁6�K6M.e�3���t��\ "��|c�@�؀�z&��0p)�j:�~Z�y4�c�ݺ��Z�)�ۯȾ�+��%�x�֯��@ 5�j@�c�&F�]������S4��x�y�U�_�fY�^zjҘ:�Ȟ8�M�����I�q= �$ק��TJ��^���*�	���O~��O qTꖃ�ŷ���r��{,�#�	+Υ�ѸI������Zu����M�N@�����x �kjus��򾑵��yD^���d����GͿ�qw\Jւ.P�wc��� ����-"�,-u2�v��X���)�ќ�49\~�N�u�=��]Z&lOu)�����V����Ȃ�31�����Οik�,��/��__���a����7}�`�>6n�����'��w�W�u�,���s����	�=���!iOn;� X���I�K�I��;\G�f�+gK�"p���"%zy����XټzY
��l�)l�y���Fȳ�����
�6��تE��L���m�~�#q@���>}�����ƠlJ@<0uH�:��ׯ���M���
g솒�a�d*Bܔ��Y��lY����Rk�k�W����r���jG� '�5�0;$˓��=]�Τ¼O�kK��Q�� ��b�p�3�3Ⱦ׮~2���D�%�ώ�G�j8V� #es�Ϲe�O|\�4�x�͵�IP����"���U"sټ��G�PenJ�Q�|��n�.N��?�jO{@�x���&��O���Q����cd��;0�#G��8��<��p�b:��}L���%D�G-p?ّJ�n=?�U�}�r����ڬl}?C*�3 "���E6��!�C">F�@W8���Jŕ8`y��c���*Chk����.^(_�3M�Ž��ɰ���I~g,�A
�a�.48f�;\�94�׸���#����T����/RB���v�]���ϫ:�ϫ�Z�:�Z`��K���2���v���pi���j�"�O�c�Gk��h(ό	>S}
uCYk�H�^������=�����s���'�B<T5��ګ�s�Xr3e0���;������|��N_���xW�Ϙ}��!:,N6].��ꖸ#5�rS��haY�X��E7���s���A��ZL�lr7;q������HBg;�B���y�%{�Q���:o/�qTO�!���ƫ�K�b�z�U**@�B�[�~}�����.3�b�QN���/�����P�<���۸�)k?�V[B&��#�<��	�VT���R����̹�A �Q�J4����{��g���;�R��tKV������ku�"�tӓ��h4=$�j+��xDװ�q�@�;]� ��M����ϒ�5�9�0q�.���΄�H4�#*��֞� ��_�^/�Q�,����D7��K����������8!�Ο�r}� ^��9��.���q�X3**��v����l�Fw]���v]���c��-
�nT�i��`�\��>(��Eɱ~m� :����1[��&�e�HF:�#d��}�]�_����gTסL�O'm^��xK��U�y�f̈�[� 6�{��󫶷�U���3�a�|�E�
��L�¡�7o'��>���OU"i*��K@o�4�����o?���4����3ϐ�Td���g�ߐ�w�ۉ������U�A,�D}�R+ K����'�gF��V���
�(S�9�t������>tR�j�+����O������S�	a�*&ض2Y�틟�T6!�`S�H�W]pn�k�N[X\�k�Z�������x�nydQ�xȑ/1�9W�tD��7��Ϟ?<�/�N�"�KYk��S����W�C6-zl�r�q�gIs����+k�[؛O�5`5B�qk�u �կ�&�D��(0o�X�����`ja�Q-]���`�&/�~ƎBNb���sB�Hl���pI؅��2����)����D��XK��n��ݦMʣ4ų�)�@��4$uV���4�1�;xo1���ln�.̾��>S��-.��t��&$�5��,�������$I�ƣ��}�vz��nь4���Q����t��B��L6F��]��m���k�#�Sl��jCUe�u����$̬vJd�-���@3��*��;�B��g����~���:J��-t�#ε��C`��AL}�:�ڝ�¿R麇�:,�⌃�ۖla�������#�ev-
n`N��� 4���3�_A�n���7��?��pF[�ģ��R�j���D�.���Y/�n���e���`ZZ���Fi�=p�?����j�����1D����;�V�$Dά �w�d�H�BJ$T�"�G���g���|��?�S|a$�G�j1^��s�	�O�	�$�&R��1ؔ:=��6�9 Y�UoUC䤮�[���<��QQ��
�~��|���_W��k%:�o&�^�W޸�p(�`K���o�����E��lR�{�]%�xR2�r5�_��>	��Š��:����:�D0��1�&h
|R8�J��ӯ'��zqp{����!;��u���#��HS��Q+y�D�ո���\J�х�%��h����w���<S�40�腎ӹ�Э�<k#
'dJ�O��(#̚��q��5I���gӂa�YQ�=I����
{_%�*����;r�
*��C��;�pNc6�n��0`6u�.8"���:���#�&�Yj`�U#f7����T,�p�����7$�i���Tuyk�,҃[_q�۳ǣ�����Q�gv0�����M�`�[���Ys8��0����eD�m!��;��5�3���`&ˉ�k�4����)h��qjx���ާm s2:^q��v���q@
�3����H�Su�?�����_�{	���)BW	�(bQٌ�С�����oB�
��e�kϴ2|-��[�}��`��C��%���[#	�K������0�+���0	��\U���>%�ZBc��G	7Jq$�;Z�o,r�BC�� ���w��PA�Vuok+o�&��Ł�v I^B�yG���r7W%1���53����#���b�W���ǋ��n�ި���ꎜ���V���'F��tX�����	�Z��°+��ň��2���l;��OX��f.�;�_#�]
���)��rɞqf^��@�q��7P�0��Em�����#��˓4��L�ZP�����-��x��6����*�'���j:a�/Y0�Br���C�2�~���Zm�� ��?�ץ7
⸂�r���6��0�~��C.e�Ee���I ��0��	��_�̦B���nO/v)�6n�B��Vp�:�+���x�_6-����i��"k g��̎]�«3f�c~:8���~� ���@�o$�劌
r 3�`xh�b����*w��B�`�M������~9׀�I
�#k�!k�ܸ���?L�xx{N;e�юѳ����v%8��D�;�-� g����X^9~q���S6�u����S(�ү�����|)��	�\���
����m��kl�p?<���q���.ƚj,�p�[Jx5�ԥ"��$�-,����E����'��KG�[a��涭<3���k8���ۂ�c��*K(��+�������w��q��v�
��:�Q�Ua吩E1/6�W��Ƒ�%������g���V����ӳ��5��X?1Q$#6���:�[���@��Q|�s���ʁ�-G ���?��[��x��R�ٳ���6ԓ/`6T����Pw�"M�~���XE��פ�/�#tF��Kף�D�Xo׍�!x���q!nT���`&[?)k�k%���o9j�G~��Q�C.����"�Tq��C�T2��ՇB���U�7�)����@�ݸL����m2�t@�d-="�,K��A�¼�Y���ߑAml���X�a�7Ou>��V���89r*�B�C��#�KU.N�4D"���I�X�G�l-&K!���'VX����R�fU��10�W�b�9�m̊��3�뤓瞦 �)n"I�����]��:k���GPDoӳ��F�@�d4�����:�؅m�ԭ�k�����iD�x��WY�tK���x5[LVrBŎxY��{d�bf�������^�J
xVu�!���k;�Ȧ)EoG�+iR�&�p)X�vzϑ����J���M�69	�w�^!6��R˫n�:uz�]Zb���I��m������6l(�nr#�����e�R N �K��K¸��)���ՋT���̟������s��9�����dc�����?��1��b����̭���W��ܫ�`�n��X�%���O�._.���ӟ`�@���ip�UL�[ϫ.<��"q�HJ�g�1���W(���{'D�ו�ŧ��K�IY�!.{�@����p�R)Tc�J$���f1��s�����q�=g��4A�Y��!l��o�)�m�ks���]l��;]���'�e^�B�G#�W��C��.v�Q��Z�I������D�\�X!ҷ=�{���E�T6��\8�Z\�5$gY[�匄�`�<��EK��w�OE{����\��8ó`z�����@U�SZ�E� ���y5-NV�u}_���`��u�UMA��
i�\��K��2/��1���a|�OZ�Y0��]�Z�Y"����G�W3��vo�|Qwg� �BB���*X��~��ME���c��f�g�4����3��t)MK�������p�P�4d�}�1X�i�:U��E�+��I��Q~	.����;���V�~���.��%�G��>v��@JAĐ�E	@��:K��"o�`(Jh��t����e:n��ua�S��B���C��܈�@�c���{�g�0WP��PaS��5 5�XX��/m \���""(�m<iy���G�'C=jz#�n��f���M���1�z�-e��~�=�Y-|�re�G?
�9�%|S�O�M����3j���2_i����Cň����5���H�5�`6�V>��@�ELǤ=��O�Ev��4=��bI�UP��K[�����EK3���8�J���Ւu��/Ғq��c�ۋ�*N�p��V��;@E�s�{X�y��y���^h�C�u�(���J�T�$�n���N�y|A�!��+�-�˾_��ͭ�ݧ���0��[������7Pp"���y�`r��]�u�mſ��/5�,5>��X ~��:�N̳�#S�:w6�B�L�M�@�3�]i��-�h)`�Yߊ��"�g� \�z�S�<I�����4�[��⍚r���_�K�
�ڍ >Ɋ��D5����|&�|�B����i^h�m���s�jF��bEܯ������!o�m��Cm�@�s���'����ԛf5W@�����@I���:q<�j�)1�l��M���}V�ӏ�����
�,�$�:��5�����7"�H��@��ua��:��k�s��E��:�[�s,��Y�92����/J��̵8��"cG;Bf��2(�>��)�g�D?)�>U��i7!%����g�w����X�qr�#�	1��au��86�ٔ���1��mcg�׆�i�+���^BJ�v�71����^�{dՂ�[�h�]@����} �t�di̦��9�g>�z�F��SL���
��ҭkSϱC*MNG_w����D=���֦�w�5d�ҷa&^5��H۔0��b,�k�g�#gҶ#�`��Ǚ��K/팒]��0�	�����R����\gP����0�C�=�IF����i�u-5t�՗ZeHɖMе��2���OӇI0_��-�Ү��Ŷ�;���ڞ|1,�9������-�g�
]�c��]�%��K-��#�1j��]8�D�8˭
�mKC���޴�������FTȡx�>��9I	r/��d
��i�W��Nl䈆��X�xH㎿������� �7��Q�m�T.P���
k�,�rޯ���,��́��l��[��M��&��b��=��~�J��X-�K	�A��^� ~KHT��5|��XE�W:�[#�E�ٹ��`ph�N7�"�7t�I�v Nj��Smb{Nk#b_�S�5S>k�����s;�$Z�f�`����	�埯��S� ��Clzƒ߻[һ\������A7.E�%�m`ߋs�:\�8������ҩ��5=��/!]��y"դmස��o�nö4/ �᪞_����c�[��o  ���jcv�79��c&��KP����_�F��D�(��F�Z;Z~à}��*:��=�-�|��4�p�At���zu�B�_���Ǔyo� ?�ȷ�,QE�I_?����[+��Ra���(�#߳T=�g�2�#��tE�/�$25v��,ۈ{�ִ�Y/dS��۾6��� N�����L)�$I��,XB��$V��[�� �L�0i/�v��Z��D�t��6Vې�%��(�@�T�g�ы��
����c�N� D��>$}�+��e�Kz�9W]�Dtգ���|sm]��u�,�Y��o�vc�ؤM�L�9Д2��!?��6��ΩF��6v��}�T�m����lC
V/d����w6�t\cf]���R'��1�3|��Qc�'T���2V����`v�xD.-��Pk�P����Kw7;� 3�J_��+��b23a��Q�5Ƞ���Ҽ�I���`����#
�(��D~��o~�w� ���/���P�{",��ق�wdv�[<(|���pUݚ�XQ��Y<{��3LSlt����|m��]{�Ү4Ѓ��}MAz��y����bHt-b��f����_�r��I{r�� ����R����ʻ���]Irb�m�w	F#)p�>B�'��0{d�f*��u��}ZM�	r����!���`ݸ_�2��^���qxLrN��,��\u��2���R��#���?
�d������ʘ;���x'nP��s��n<ד������	J�ε.���(���h���V��9<��m�K�cVC��%�
�0�j~��`�l�xQ�b�s���v,���XA����r�g@��h�:4��x"lG�X� ���դe\�߂�?����>��F�=�)ԩQ�ڝ?�O�S�#�Y֥�1�^��O*��1.Ⱥ���̀�?��E����^��`�io�q�����G�_ Or�VHm����
�@/�?�<��-���2�O�=±��Kp�gP�X4���P1=
s�IIؼ,,3j��`z7�.*��Ξ^��L��>4���9��y&�f���$���p�x����ͼUx��9�䌬��q�[��-�Ýے�K������`/%� �-�s䃃�<C�cr¯ƽ]&�V���)�M�+d�(�sG��*�����Yi��"+�|g�;ۅ	c�pU
�ʖ:��_�|'a�����?�_�Z �X������+�2��W��]�)�2{@Re�&*��?1�XN���5wu����XLɘ�ifx�%��7U��}B�&���bn��Mؠ��PY9��@��T��9�JO�_��r�jl>r��A��v(k�m��V��Է�ʝi�@�Z*�NDW]ԭ=]��hl�ھL�USO�T�b�L�6���ؙ�!SD��?s������|Lv��7�/UЦy5���V)�8�8��生��\&-�d�)�r;�V�qޗ�i@�AfZôsӅ�T�(��u��c������z*f {Ʈ(�GA���&�[�=�`�J�R/0�T��@�����8�|��w��L3��L����b�} ���=���J�f���Vǋ~�X���7�ź*̈�n�"Wv�ok�<�E�p���6��x!�Aɣ����ߙ���	F/a#4�ObV�,��ۑ��W�T�+�0U��1������N���q�1�[�ȇ�>�^��!b�6�o�0 {��,=�N�r�מT)x�;W�dĆ �i����u����}��}c�A�%���˟��ح�L��L�`=�/��|}�'�g�W�m���'@��-��xHѪM��6�u��cbؓ溪�)�	�8i�o�/�]~@��W��5�"�%�RՒ���ѦE(++H�WCE*��R~&��~5�h�S+�z�ԍ�Ce�*��
T1�E1�t��>��,4[�az$>�7�/c�d�����M\�OvRvA��ce�y�U��{%�ڋ�A�\-q�ZR��8�z(�4 �L+�Hn�Lv�R����!��N�MH��b3�)T������q�q�%z�sװ�Yy6���v��W���Z{i�G!�<?�a$B�"�fM�N�!%!���X�ʎ��^�E�|
���6ÙJe���25�Ph�俲�����<���	d���7<vo:��9ܷ�@���ށږ ����Ewr#�V��~�^����_7f�M{52L�bvE�����`y��������얔һ#Ж�ӯ+����I�}�[��V�J�H�P*�)�_MCG��lp!���[ДL��x�$����nr���B`�^��u��ͷ�c�'Q��9��[�lqW��+5~tY�00�u��*�pD�Q�Ly�h�T^��8:�b�ZK5�U��潠�e�`Q��."�|K���,t!�:�nh�v�`�A�F�!-�>����;56Q�֕�0���U�^����4�_Zb�A3��]�6m�\�䯣DD[�2,
��Ō9���$V(Cv^�0�|��7����L�ъ�%��9��I�����k����9Q��~Z��|��G����|�lD$
Y�d(k-9�ɘz�幧�U�_{U3��\=�]�u/�|�ǎ&�❡3I�=B1 �Z�229fA����#���%/����{��C�X5)©4=iG �h�3�OX$)7pqQ�;���`]{�J=���Y6�e��Q-n�K�5o{�m��[�Z3eF�Ϧ�͇��"�l��8���1P&�G��=�o���	3L.
��F���Ɠ��_j��8NDi��U~��]%�S���*�O�Y�ޖ�T�r.���S�k���h���iB����%z0�BVMvJ�Ms>��2>
�h�8�^/�����^�K��������QJ��Z�B4�0J:2�Ua�Š������i8E�k��5�s��d�*$k�x�^��7�ȍc?��"͋R����eI�1t��	О������"�ߴWb��i:(U��~oA$�:�z	T�POJ����YjQ|7+��M���E�<��Sp%9�+cn�d��u�.\4��1N���?�^"�Eߙ��a�,�Yn�/.�$�$��#o8���
_�eU������Y��Q��Άr�C��UPc����	W[�u��<��7��ָ Id�p�"u�$�Y��zҗ[�%N	[�bɬy4�QN����~�CK1&�|j�+�Q��H2�[���m0vgE��C&�k͚JC���S��{3�Ƣ�J���U���4�i�v80�=��/��]R[���X� �nц=��g\��u�D܈��FZ͵�=�oAkK�0� �r�HĞx����)�kB��1E"]��o��D����������hix@�ӭ���W�[�{N=�&��<QgS�Ѻ�s��JcjG��M���~��,!��v)�I���-���}j�:�(��"Ia�\a5V�۰�9��ܩ��e#`�'���NpV�Pe�Wz��L.����T�B�|9��Z���"��S����c�Om&�0qvi�8������Q��m��=�>.5}�%�_�BA�%;��I���F&	���~.`]*GZ� V�xY��-���q�#/��W�:�nP����)�t�+�.tFQw��r2Z�m� �����eOH!�����/�q�<^2� ����v�"��4 ������)G��s��ǿD���!���n���u)���JS������&���6_e�G1#L��їG�}���9��ߝ"s��,����r�͎I\�ʁ*�M=1C#���jAɕdW�.�?�Y�o�f0�J��Q����O}~�V+�!��1i��jdNmG嵤�.?�Nǅ�	���,*z�E�>�֒#T�8t��T3�P&�� �9����P�� �8q��}�f8we�k������VAEP��S�W����Vb���8���8��:|m���UoqX5�����c����~��h̓�@���>���{̭�n��s	0#	s�ER�_N=��U(:#LJ\hϿ�T�,<����zb�*+�F�T���Ql�Q��S�ݳT/E-Du�MdXE��R���H�]��ي?%�q�'�f�u&�����R��bt	��Z��!S	~sI�V|���\�Y�� l������3S�4�W�Z1�b�o�*S���q摯�s} �I2۬��l���=[�F�E���ď+����Z[��<WzS�����/�#S����?Y��O�*�X�D�b���%�~�5Zu�H��U�R�(��D���N8�x��Q�AD(&5��]�����[۞?,B�/��C�~��L�M&�XK��ى�'�K�e6��3yVu��%tq��a�<��w�8լ�3�#��.��_h�mgm.���M��Y/X|EU�c�^sr���qf���K3rfG��S!`8wj�S���7p!�&�š�����	��5�P��CH���(*Q��[XoP�C�G�՞/��W����sFm=ġWIlv�"�jŉ�g�ImH��x}���\*���P��&��*#�we�����)�r������`�@�~V�q���R�R�H�=hP���~-ۏ.~�4�e�|��P���:r�����v��CQ�J��L��=�'"����y8�p�Pt���ݘ�?��~�iKq��qd
�bʅ��SC����a�	���Q��l��Ƥnܥ��e�����= �p/�	yHl��j�06E�dW/+��l�����*�T?���4+��g����#j̬�tg�Ԁ�)}IY��B/��yb溎F�K��[� 2(�5Szİ�����0c���s�o���
��H�*��۹�2��	��c�g�JL���&�5V6�^�}˽�~(�(e��"�o�����YGa��C�tܿb���,�,���$�����;�+��>oՀ�3�"�e'��Ʀ��)@=�YJ�%@�PJ��G�X�C8L�?����to�N���P���������؆nL�� �845�mk}�O�����[l����IHLIuG$�c��d���U�&u
�Z0��1Ē��qB��sR/0��q��W�����o���)��A����Crv�"�#�:[d��:2������it���BR����pwm]�V��MpB� �V��*��~(���O��Bb���fŋ�"Y.���Z��^a+{]��ᑩ挸.-��%i���;O�X5��n�`��k��v����Z2fv=������.-w���l'���W���;ٴN�\�Y��K?s��>b`����E/o���`8|�sΞg�bOm��}��g��!GFZzU�֚VU�;���4�$@i��T'J�(s�2�C�p]}��~	mV�u���?_�S��=*��w��ç�,9�HB���j՜���l��򌁜cwY����޽rr��p�R�I���hN�W��al�kqA�g�1\�ХV�!_��<��-?���
�Ы0ٴz��E|4~�.��~�a�{�;�V"Y��@SI����kp'+������<�썄B㧊�%kVk ���@ ��_��E�M�t������l�d�b\g�)Z���{���q�!���n�VS���Wx�A
�D0��ܫZ�A������R�����) �l�ؘdL4�ь�����㶨\���Aq�����b�
�A�6�ҕ/�"fS�q���4t���a6}��w�OvI��Ա�A4B�̪��������&������_b�+~R�m9�zC�*��k5Ŧ&xцT6�!�;٫`��:�Ξ-2`�R���%X`6���=�Sx�pg/@��P]��˷�|�%�K�W�֕R�ve$,�������Va�;`�K���#;G���Vz�i���͂ݗ��@G�J�ERH�V��}�����\��M]�?6�@dY�W�b�ߝ=��G:��U<U|�ٻIg��k�u�A�A9���j��$�x3U�/'�-����Ih�#��s��nl'���Á��J�8#I��I��F���&#�qR��gX����
?�V0��ƛ]D�0ź[H7Y��7p*���]�j�͂�h�����2�����V�g���~gNj��7ho���+W�W6����Y'34�5�rU��&b�
\;�8`�W���u_���#.����U�?�D�2�N"a�x3P�ut3 �j`�i�e�
�sOb{N0�@�"���V[�`Q|Z!�"�����y����P�щcqM�&�JM���@��a���?���qO���@(�W�Wo��;Х0���o���TЫU6�ȵ������8(��W�Yx�X���i{�d9�.��*��}�!��O�R"�1��Y$�Mu5{�&9��H���X�@wvl�������9~��䡐L`���rڞ��9/936�fjQ?8yP9}e��9z<�/���>^�ʛc�7��qklD�9�p�aK�M��&|�1�1�֯���O4����i[�!�IIg���������ߨ�S����b,���V���>
��������1���K����|�u��fV�#��##���)c3��`�y�Rښ��o��M���e�pJh��v�� e�m�JoQj�d�P
0ZC����4����[�0&�7����^���' �\xI�x�j0xF��P��O~��2�b�F��4�B;�Y �
�<��Ʉ�t�VtF�B8�dl�l3�Igz��p���(H�*�#n@%
*�@ֿ��q����>>�� ET��Hg�g޾�*!$����T��l���iG����M�:/���t��u� d����k��o�U�(�w��|��i�K�j��J�X�fD:r��1�ڱ�ڀ
ui�r���6���R��� ��]c*g���3�K�" ���T��Ay�L���#�ـ94�X�K��`�Kldy�x�W�@wn愤�Xt'넺�!�;J�[�R��7�X+�������2=�(�J����n�܋Ï6�8�nu��t*�C?˃%D�����e�&�,~��-ra}��v��������pS�'(��()�q�_|�=���紱���OF��&�".�9�a��=��_� ҜG�Y���;W���s߄�n�s��3�gS�%/Ko���#>ؼ�I��F�\�'�iem�,;/�.��7"��m�qžv�Z.�@�`����ͣ�\1�1����/\,pNC~$���"��3�)�pӭ�4ӊ�|C
��'`fz=��_@w�N�c7[ժc�������up�<qD�_���I����q���GI��Ts�"a/�����Bp-�]#��vD��s��U�~u\�E�T8ߎ|�KW���f)��0P�ܯ!�s[FP9u����~��qد�;����UАQÚ$J�:5��+ܗ���f�r�9LǪ�tŪ��@y����@��1�
�%��;�KBD�9#�z�c�崗U�Z~C����!�[Ή��ld��1�T	,���,*7�}(�#�,�S��F�B�ȯ|�5��y� �&�tPF>~ᲈ,C^~��ܛ+S
�o� ���NȖ	�݌$u��PH����5ʬ����&IZ�_-M[+��"��h��h����p�����k�U�x��j<en�GS闠F���
��:��?Y�KJ���W��e�\[�]pN��˔C�wK5�o�2���T�'�bߘ�m��~�BW2�+)�۲];$<��-.�� = ��4'��5T�.��<�!�Ukp�;�C�|.��g$��������ɫ=E��p��6o��+{F�)]����H�N��Z�O����V%��n_���Կ�OT�KQ�MѼ�<��St���b���⦮�:n'�Y��V,��K����
�FS4`�������i�z^��!���|B+�Or�;��c&�B�[���W7f�-} ^�����F�C�%a5�G'Q�f�9�b�X�jE	���J��6Pj�m[�"P|�E�p_slEiyR���m�A�O����T�)^lo����^2R66���L���}�9o���B�N�[qF�`���XE=��zap�� �W��C�6�0��롄؝_gc��x���S��P.?L��Lu(���ײ������|�L�tm����T�v����\Ua����?���cx��+�R;v<�bP\³18�y�b|�|���1<�ƾ��Ϟ��i*w��W�U~�Ǯ�Wv�}1�y*�b&k> �-A��V84�?�(��(3��oM�0I��k�з	���1���� 
{E`�|��� <$c[t�����|�i����~��Q��p�q�B�ln�nZчP�1�9;��~&,8�(Nk�H�a�P�,}&�3��-��F�3�S�Q�~�����2�B�ذ�u��S�F�gr�h�r��8�}���,i]������	�u����-�m����5�Tz1��N��uy�o\�#c�Pt����.�w��=�1O��u5��p~�^Z�������٩G�~�׀@�
�PY'A� D���w��� ��������vPT4�ƹd�k)�k�(��:3%��@�"[�D������8�e��:�p�M�ӆ�����_�پHPʦ��v)&VK	�I ��+�C�����aԵ����G�/w�:�YKz>BՃD<,�0�/FH�o:l�s��ECsJ1�e~K�Q���ĺ�8�Dy��I�2XZ���O:�B|��il��~U4
A����=���uM۵�s0���K-F���D,�5h�ӫ�On��[q0&Ui���A�]�����I	Wb���?�s[�.��bQ ��˭b�^�萖X����F��ء�68�.�T=�$��Ǘ��N=��`E��Yo2@@��������:����}!�{$9�ovd^��U�Mĥ4�ﳌ����":ŕa�a�l�e^�ٟ����_�v~��5'�nD�:q�*dj��|�pt�^]��Wf�ҵ^�ѢǗؗ�"8���kT���04��j�j�}�rބ�T��t1�7�5�BL��]T��rn��#�zV�����6�Ӕ��$�m���}(�c�O���"�AՕ��(�H@q�F�f�1��(F&٬L�|��Ch��6�B �Hc�N n�]�v�f�0GV���g�Q-p`�_��*�S�<��(��J���x�ۖ� ]�����~�	P
�'��XL.ӌq�{���aj���B���*�R��Qc1D��3y�_�̅Q`�}��_�=BV %Y݃_5G +�WD9��@a�f� �;8D����Tn���}7��~�i������D��?��:z��a����;�T�AVMK�G��d&��f3�c�6Vz���{��8V�$�Ue�f�u���?��hV�6�Tiޥ�K�A8ᐺ(�S�#��8�P �c����9��$�k86F���X�H�/�p��@�ə��Xǥ�ٷ�#�:L?K��ߴ����@�d�'�W�p�)���>b�iJkJg�@:��[Qx�(�n�-�W$</>K�:&t�/�IM�_Uy"�:i��jm�k��"cmQ��XZGq���Z��;�w�š���T�0�Lg�����-�[�n~�_U$�Ĝ��Ŵ�g�x��67�3�GH�4�6;�=|�\�Gj�e���-��fx��FХ�0<%^�0R���5��G�K1�ة`Q4�[�G��r�P� ]�fҠ�N(]���Ѣ��86a(P�"^�cpZ��D�
@n�#�z��i��J>;�w'�L����È������^@96(93n˪١��1�U�m.��P3�r"�*��2"�����\���S�U약����t��p�3��s��TIk�*��C�_���'&}���%���h,��g*U�;ެ�ZQ���O�Rs�\�s,�9!c]hM��:u7C�D�{����_��gξ<0����ZdRX rŚ&��XJ����g0��w����W�ۗqm��.z��/�-���t�F��ڿ�5���Ja�3%�s%[Θz�z�S�>�C�O�6����c� <�����J���`�P[��u ���#�i�n'���G�6I�%��Y|����\Þ)lr�wFvNT�â�"4{��'(�'�⧇Q�m�h��e'o�-���+�:
�)0qQ}@�|�:B��ƃ�tM�褚:g��}4N�X�)@��{	��:���\�?PZ��;�G��H�b��e
{��4��3[����`�c�� �3�t���lgtgҪ��J:�L���b��⒀���9Bvꕗ;���6fJ�#/o�T<f�V$v���,&3J����&-P��|;�;W(ҳU����^F2Di�?i@�
fgX++�'$?$��]R{�*�02z�Kh�֬h�,$U���GLd�����覜��.F�/e��+8`�>���$S_6J���4"[ BDָ����3��`o6��3j��b7�V+&=Ns��H�Y�)���S����3S��lr��j*�'������y��<a2�}������H����S3m\�av�B�h�=&��<yL�.�:�{r�n��_dГQ2�[�|k��U�܎�Eady���/b�����\�X_��h�Q3Y���5��a�L�+���^��3�T\���@��ͯ��]O'�('p;�q�K;_��Hj+Q&]�y�xF=tl�µ\v�,G���(��3t���f�r���@��.[���o�W�$���.}��k�ZIw��B�rV��E�,�7�H���|�	�}��f2]��ш�7MU���<m��!����_5N� ��r��J��؎4�Y`�ôo�c���/�Z�\�p�0 T.�%*�8#�:b ���ٌ���6�0��)�k���]D� ��v�-c�p/*d�#D�D�/�)�ЎBW4;1Te#���V������̪؛���2P�\�(I*ז|��S��V� t��A�%����+<BfaO��\�2J/�7�H��İ��+�s�;�6.O)n1������I:1`���tQ���߼��C��r�2Q�v6���$�����U�GEF�2�H�����g!a��!�N��-��q�/;Êe<�=L�7�R��dcR�
@���F�����oQog��v�K�W>.�_<G��U��rg�f�N�F�=�	����S���Q��ڡ��-�����)4��y k��,6 V_��Ӷ ׻��|Ċ@N�!��$�ʙT��XU��!J��A"���?�a��!����F�n���2��ʌ��X�!��a���Ru�1������l�?A~����;W��G���n#�ø�C�0�&~��]������ؑ�t��vm ݯBfjD<�ŃiM=��I�A1���(���X	Ȁ��0�5��S���c6�S��Ҋ��v��!���<���}c��âs!�}=��)G�N��}S��U�Bt܌���VeB��}lH換I�Mj;^�h���)_�پ9_��s%0�g<u}�3�g:2u��Η_��О �W'Go�zsر���}W�K}|�imv!b�h*�;��̐+`������QC�<՘<�@���oW��Y*���c�Ff���(����!~U��q˴��U�����}s=��Z��`�J��� T��4�Ӌ�5h���`^�(����t7!�G�����m+�Y���b
��T�/�3�ͺn�����C�l<z��5
z�}��l�n�='o�CZ����5P�}��{`�0��f�\CN� 5���4R��)k����>_<���i�B�m@G;�x#P��9���M�1Ģ0�K0�i�&@���+?|H��9*;:�?K����M�H\3�����J�Wy�f��7�7���ݛ�8/��g#���؝�M�Շ��zB6I�3X�ňuB�(�_��8�oFm=��kz�����)�"��*[�h�m6��0�Ze�]��3SFrc��L�GAD�.���U�l���.Cs��]�� ��e���MQ,��4B����.��}/6A�h��f�_�B#F E�x��<�����e���˪�_yt�%s�b@�rse�mV,��Y�^���`r�����T�QB5-q-��X�D��!�r��Rg� ���䭸7��.�}�5�	��ﳢ3�Q���=���
T�!ţ�˾���Se��[P�Plx�iر|�ڥ9���s}S�8֮L<&k��W�&|B�V�ܭy>����|#:v<����i}�]h�+��[�ޱ��*�q�0��;7&i��:q���į��vN3-؋U_ϸ��8ǚ�C����wv�[�)Ö�$����I��$�a�h�Y�2d��D�Ҽ�]Jp�I��71��;(������bm1��ZT��_��wݒ~;[E��;��sݘ�?�!B�l1�̛fTXӯY�t�a+�9��ՠ���w���Q�m��緄��N��P��X��*� �GN/JB#}���dR�]�v@P��%rC�K��e�t�{*տ[�I�@|���*��c�G�pL;���U�-��n�D���	��N��j�y�E���?�t���=��b���8JR�%�z'*�3	*MA�)c9��%L�kh�#QV����Ppp�C^\��a��I��gC��cE���]��͕�)�Xi�e�eC��a�Su�*Q_��r�`9Ǻ�֑��I����.
_���cJ1�,}e��{�T�r��;��9k���i���i1�)=�G�| ���a���Dy�՝;�r�G~�;�Tn�ɀuY�>�N�~���\�#�Ƣ��D-�ʱ婞��}�!���=��h�>l�Ӱ�SP�G�!%�(������ن��~��C�{M�F��Ü,u���B\����s���LM�+1��p���H�46��$�����֕�_��{OZ�i6o�nv,"(��Y���/�7g���2���4��
��(�|��5���L��z��pWlR��r�ɤZ����P��"L�1��c�1�K���֣�hFdLZ<!Z�\:�Q�SS����eĭ�1U�!��G����&�j�ǡ��~�"�A�&l�
�_�F�"��ÒT
��!6���@����ф;S�|GE"�$���k�:����J����s�A��v%z�,y%df�1O"x�c*Y��7�M+ydbs�紜ɭwN_%����v���'��k>	r�n��h(��	Ԃ{[�Du�j��
��m0�N�b���xa��6/�ٞЄ\�w�Lw�ͽS6,vG�]��x\�]
�xq�'��2�dH�˭�oZ5���˶8�A1b`�H �~(/�#�9e ����t�5�ѫED�lRs^����Rt�qOWa<}��߼C��9͂ �u�#�����M���>������e��}��c��މ��UbN��Z�wS%�#A�OpmD?���q*��3��!֒�y��[ B
�)-ǘ�I�J��;�Dک��b��*[L5�9��A����Fq��);���8�rB2CXbu<�Ng�(6���U�87be�K+�,�P~ypF���>4�nW��/l�.��Xs(�H5�o��(���*D闎R|�U>�B��&��4��U� �a/GE�Z��}��"�~�s��Fq+�6�A���Jƀ&~x(1&P<�����ˡg�����bh��eW��&��Pg>��
����[j_�u`�0Z\}s�d�Y�t x���O�Y���u�^]2��(/�3�J�D�eNg��A������f�fW�����N)�C��m����#�0�%��3�z�[�˛��j��fBZ��f
�҅T0uaA�vD��z��4�t��R���O�|��1���H�����MƄ�:�Y�Pr�f.Ō�������%<$#/�g�<�R�\��!=���U�ɴor���Ɓ����J��g=;M	��QD���|�AI}N��X��6��~�J�8$�ſ
U��B"I{(��#�$-=������+��d��$mi�T�����j1��ɞ����Ľ�Ó`�ȣZ;���GV�E�E�n�p�x��AtWm*��:Q9�#*���)xR-��rR��0 ș{Y�B_�~���'��^uF��&S��(ؠ�91�9�E�;�:��_?t�tq�p�
i����6�¹s��b��X
���o���UƸ�ȅo�4�5�|.>-<�{��H������G��O����\f��A����#�~�#���~mqo����m�1��5�JCt����@��!�v��p�	���()���]mR����k~qL���U�X|�n��&����ԡ�Bt�J	����$����Y#y�'�����%��L��f3�M7*��[�;܅�4D��5���L|��7�ٳCRd4�[z+q"��5�έH� 'Յu�QH�����$!�SZ4����R	A�s��C�c\/���G��2��\`�0�I-���xQ�[A�[uA53.��f%�FV�X�?��V`sRf�����rz���xB
A��h�ѻ�m=x��(�������7�i�j�7���m�KG�+~�W�y����G��?`��q%�ϓ%Ɯ8������Ǖ��R̂j��]m�Dd6���I�1��MI8lT��V 8'?�sn԰���,���LO��T��[�*�K.ݖuӒ���u��̵�]ZKa6򬄸�ؓ��ZzO{Vv�u-Y�#�xʫ��y=�&�,������A��oR�0QǛH[��8��%��Uu���6YM�^��k
�q���$�(:2��~OJ_(�r��_r^^aJT���VÛ����J��mc3۠�@�ۿE�h�XcQ�B�A�9�To�C����$����q�!�6����#�0ֽ�հ���Z+� j����i�y�-i�q�d���W\*}�O�Fe"tl�V/dQB���>@�m��O�OI�Ky���xS��DH-TΊ�	�f1!j�q)�&=��\e���1��� ��s�|�.ra
Ŵ��3,S�|�������/(W��O�~�2�_o�%U�K�P���w/�I]a����*P�L��ď?��3�܍�v���K��Y#1�[���Q����'6���7��p`�^�#�Z�Rv��?�+��4��@DP�D5q_a�<v\O�ky�b|qT����>��y[�Yr�.ŗ����GU��kh[Y �m98��	p��k���yn`i+�{��K�#]�e�ݦgU�ۅ���`�.�PRZ{ițbڞ�ҳ�b "JF	k��>V��&s�����j�1
�r"�W��@�cj�K��U�vQ�XSƃ�ϙ����y[N��Pu�V�=��{W	�ڇZ�d�uQF�f�v���K3�����^�i�vɋ��b�-$���Ƭ�:DGN����:˙6tc8�Mu�k>S8H��U`���^�e�5�pJ+>��^�O?i�Tp.���.���%*�N81��gA��E��,^���Ɖ�=_eF���?#�s2��OmXq���	X�u۬�$����ߥR��~{�sc$඀�L�.f����-[��]a�0���t��x�9ܺt��{�MN�p&�=����ɵEZ�I4��#!�a�gj5��,[}�r�"�f�쇬�j]��4�Q&[�g&_�W�0%7@�E�{�xه`������,� �Ζ?c��!��pR^p^8���,�[AqM,�X��,i�a=D�5��y�3R��JЈ�b��T���_P������r��X=~"&�L�x�sB�ҧ�$��&�OH�Z��Heh`k��Ub�`5�7 VN���������>B��Xf6ؔ��r$-L4:|c��3u�V�� �~E
���.��)��[}��~eaF^���縵����S�'�~�/4aH\_3���+�үˠ멓���9r�R)d 萀�"�g���~��d�n�aN���@����+J:s�˗�Du��2gZ.F�֟q�?�gm ���"�_L��n �y;jh�?�D��B�[��<�}ɩ턣T1]�G�A�Ih����n�=�9}ӭ8�{�{��d�;� g�S�F3/Zy�=���[}��\OP����5�2-�㐞�y"�e{Q�ϟU�4IwD�`���� :��\Z/� !���?�Ӂ �Y���z�ׁ����VQ8�#-_���t�a{NǤ�t��:&�}t�gp�pPrˣ (����0�T8N�ok,�kG��~�<<e��_�p��9�� �I�T����U+�����h�ɑ��?����=���~ ��	LS�=�����Z�=�fl=(P�9r��"�$X����|2s-4x}��R��������u1�^ T�z�@�̄�Y�{�N������f]C>�zOe.��|��� ��b�$�Hݽ�s?;P9��tc��B�9&m$ʹ���1.��V��9z�B)?|8�0Z���5V˜��Z�;Q��,I+Wo�T~�����-�q����,��?W�B��I/�F?�k�)Um$�0�Ř��[�]/Kvy��/���%چ�[~��t���5Tp���#pw�?�.y���88�f���U싧�0j����|�I���b��G��ˈ ne�ܡ� G�l:�|��2�>(����2I�3ǆAnB飡A
������3"y(�9�,�bI;4��[g���&�Y��ύ+(���-��֬����G�����d�I����X��������~�8P�ty5�B��^����i�ʃFG1�H�����UR������J����91p��%~Ӯ�*�]��C��� �}�|�	���G�}�"e���I�<N���
ČW>�6M 
krJ�6�m[�D)j��<d�n��xq�c�O~�+|���3ʼ(㴛��ÒD7	x,�-7
�L��>�B�`2��#�:X��\8�5-��붚��5_� Ј�]�=$5?&Yyvu��f��PqZ�|�/��G��rO<}�O�����ꏿ�,h� uQ�WB�]Ai����}( �x���$�:��:&�L?s�o���@�����L"!����XU�(Q��@dX��X�a�z���o`)�r�u�E,wx�\/�p��Z� �#{��*�=ꑸ6AbV$Ɓ
�UC��T�|h~�� ѦP9oCe��&$�'#��T����k��@�j�³�rJ!�&	�%$"��36�M����\%3>���ZI���;.���ɂoP^(T;�����
`hʷO���d5�=�*��1�����r�m�˨g���b���ړ�Wq�=�NV*֏�����$D$�l8��d�?�s����
��UY}�G?ҧ`=aȔw�����Ak2be�l.�4��Q�	6��lCLǈ� �Q|��S�?��0n0������-�jL �<�l@m!>1�+"�}Zpx/ +�h��/�3�͜�?�pz�����n_��.�Nر�Z���#���&���z����� !�S��YG��n��Z��(����cw%�N�=��n��'��.էŎq����4���ޜNf@��Ӂ_�ܫ%����l�\c�9����o8��9���؊����4��w��o�'��n�ƺ�j�\����0�!�{�(���n��o,�*W�o��k1%p�@ͣ�"���˳�Tn�t��$��ch�b�^�+q��V�ɒ��*·\0���q-z�Q�>l\�r/�� 1�?9(5��	
�/G,3+:a�-�3'E{7�btS���;��1��nwcH��pSt���wN	��RU@S/�=�E����$��\f,X6Z�hj��g�����<(��[`��o�w�e"y���3$��ةb����)��6e�3,V��� ��<<����
�P��\�c�x3p!�>>����Dvr8Hamx��ӵ����~��͈��-0֥Obc��<T<�S7kC`�1ۤy��2]s���/�wG��g�_���L�g!�����������qk@���Ī�y�x]-(g\A�ԃ����������ڸ��� SJ��$s��Յug\�lc yB�TG~��tڈ��t�fYa]+�%�����H2_�.��M	BzIox2h%���D�p��X�G�^x&���۾�mf�rS��#�Z�O$��Y*	��Sy�w���_8��s����gOm�M#��wep�r�̆����,E@$ y�M(䥝��p�f�;�~1�£ꏢSH���Ÿ�e�ޱ.�ל�fU�D[h������&�.���Y9�T����d�o3��ԩ\4�+"��D�J3��?Bڈ�����pT�MwD&����n�od��[��
5�t7#�����c���O	��Ŀ����%_R����u8���ޤ�����w�ݑ��#އO�y<�~�<���;Y�P��B@�C��t8�+��R���|��:�W
_~/�cgNĒފ8M��9�M傅N
���*�#L/E��Q3��葋�;u�%g�Z�8����Ė_�qA�����	0���Q�����}2���+��O�)��ׇ_�ܔ�
�sK)��b��1H�$hc�!F�;S�S>�-�)��yI50�P���:B#���k������]V�7��d���>x�=����+8�h�ꄬ;�f݇(��S�I��bpP2�ѣ	�kߺf�@�ݺj[�A�M��O5.�%��+N����B���֘��G�y����\~Ff��x(fN�U�hP+FWƭ��Ys�_�H�Fn�"d�O�X��h�{Z��Z;[���
��.�RK�g�ybEW������<�W���������R*�N���� �����_�6�o���l�O\�L0��>�������)<\�]����\e�q��Zq��w�fn��\�σfLg���i���y��6^Ltb��Xi�D6���)��3�9y�>pGʝf������:��!��8�s-�h㇝Oύ��ƍD�CKDw��.͹����)��N���:lgW;E���&�7)x��\��"���ݳ6銞ٍ�#f+0R�z�jM�K�
���� Nv��ٲ��b�zv�d�:o����	@TF��3�,{쎅}q�K�L n)�?~�w�9�U��-���ɤ�D��F�U�Z&W�ŕ�e�w��-}�i���:�w�la	_���h�������@�0\��c @�Wd2×b�c�뢮� ��0�j�s������ +��c���@�-YeGf���Ù��� �C�c�0��̼#Ke$c��"�>2vѼm3f����W���o�����kl�d���Eǂy��`�THX(] �fkQ��9F�_�� ��m'��6���7à���?'��n���j��@X�*�;Z�p޷ZU�3����A��I��"��ٗmC��[�n�1{�V�`:m�Gc	�������I
|a?�z��=kƠ��0�ňd-҆�k{:��v��^�&�&tJ�XJ1:i���4wX���5I&�Ѭb��`d��,�>A#&YI�L���|[/�>8�1��f^�r>ۮ��7IHȩ\�[@Ȱ��<����p1X��x@F�g�g�ԑ8m���ɫ%�zn��7��n����<U]-�C��
��#lh��#�k�F�Dg����NP�1�Y˿D���;ݬ7s�|"�6���2[��(�/PSE���n̦;��1F#��s�]Q�{���[���;/_ }7%�L�����p�0D�I�4��Nr�SJ��C�gޫ�4����E���ه�d��ܑ���0�ݦ��Y�U=ꌌ���d�g|],T�� ����/����.��:3ņdF��>�od��h�C���b? �x�eʬ�|��0e����@Ց�o�f9�	}�������yEd4��ZgE���Hi����G4����>F�7rD��E� �mOm��k�=٠LR�/%�g	�xЩ_�n�?�	`�\��x>�"qs��3�\Y`����1�a0�����s=��^[�JOu-�<�JH��	$(h�j��>�:R�0ߗ	�]�XCBJ=1�VI4@*��K��R#����I_ż�<,������N�x�b�����G��َ�~��s7%� �=�d�!G�3����l}^��;ƽ��&Տ^Q��y������8M�;2\� �2��	+Z�Q$����+ɳ�yz0�Z�ƈ�cmB�g_��3���X��f'0�0kBs����%�~�|����dڂ+y��Nx�l��xM`*7��d=z<	d��wlgʍ� %5����5���qRy_���:V$��a1�
gM�Et�B�Ӵ>c>;��}�����PՕq���^�!�w>���Ԗ�¾��w��{�@4?���ak�/��,�J'���M<�� �@�X����jw�����n�gR^;E�e�k"��77B5�H�xP�Qzȫ3���q�WY����a�<P󜖃L��8�Q�ӵ�?�B���T����vM>�ŪZP�
��r�Q�,Nߚ�)f�  �R���5�x����R��ڃhP���t�U��d�? �������\{޼���Xϰ\P8��*t{�����ó��A�E��$����\`>��.�^�T]��F0ڄ�y/��y`X�6 o��Wbcɩ�3(>��Er��![R�����rvq�<���y{mo�ey��xތ�=*Nv�e�3����R"��ϦQ?�J95c��u%�^���V�pj�_��OiOn��}.��@��ضK,ߪ����.���Ғs��#nqZ1���מ�_����KJc 
��E�	���q������XQa+�J*	t��k'��7c%�{�����'�H�S~�Bۭ�~<"����y�{�Q�d�,i�b�*�$��ǟ���_�v���i]*bK'8�%0�ь��^��i�=���ȷ\��ȟ��t����j5����G��:ed�NK�S��<�e�mC-C�t��,n�.�6�k��*˿k�tU�����r��YA�UY�3RL�x'$2�����Lϣe6Y�g���!ŵ8BJ�*|K��7/sEmD�N�Om)3~�������g����d���JV�<'%G=[�EY��@(�X"j��I���t=OH�f�Pj5�L�L-�0���#XG;��]����/�Y�mp�l�-� 7!|���y$�xgtO῎��ˉ6��sh��b�&ƴ�+?��CI{���$���[�<�M��7��0x��~��	���V�h �O+�)�Ed���8+_�F��o:��{"4,�<FH	��rt���D������J0��\�G�Yᓰg p>�/4����|`x#P ���MC�f#=���N�}�j;"F�D&�i�&�_��E ��p�ߊwf�H��4�@J�"��"�[���lN�ٙaH���ñ$�x:ƞl���� LL;�~�`-����m��ʍ�ͱ�iFY��$�bYߵ�,���X���7F�GIת��6�Wy�?�ѻ3ʘN?�����^6�3���h���ͧ*�ߗ��en6H��)���x��"����1�f�wJ�wi�0P����u�
���j{�,q�u&h�P8���M�z���|3�I5� ��N]���ۨ����u��~iҎL�֢\zY%�_��j<X腔6���|�u�#�;�6�̀�l�,{���wZ-��$�����KĹ2.,"����+G���Dk2��-����Ϝ��9߀� �c�}��ݻZ���ĝl=C��ryoG�J�xƗ����y��."��ྯ,�YL:r����t����?�=�r�5 �4��3,��9�cS����NG$0%w��c��޳AO7b�(�a��:R��}��b�@���3:	��F�,O �,��m��R�ޔx���& 8��2u��Epy�k酞(�c]�i���R�2,*����I�˧�_�׶�aZ�aR`K�K��\T��y��^4���y�g4k�{��~m� p��_�KҮ�����w`[���3���{o=Ĺ�M�yq�D��+۹�>��q^07�rd�98`��|&��8]�E���M��C*��Kb����]���f@y[w�Q��G��(�M�g\�"p�6 AH���5��x]U�7��|n�[��"�	�9N	��0�
�Ē�kTY1���xT6hҝ������M�7 �!�6%��n�|�[�T`�����J>$v�Ȋ��kx���n.��xʌ�?��f2m
�5�~�+NZ����[��}B�@��ǲ��B.`���X�1�cBM�T�����桔Bl�W��bČΊMt�Ӱ�|=��q3�9�.�D4�ր'8Y?%�n����n�b=�
��X�9��"��*�+%s�V�7�p�!��WAC���0�)�f�U��a�8bfu�դ��|�j��MS�,A%ǣ6�7A��$y)[m,�:�HqY����6�C����3r�`�q\���v�E�LhJI���WS�P����Mi�}Ww��:�~Pr�oD���Qf���A;����-����r��xP����c��g� �;�������ײ���|�+nLc�g��5�L�号0����jm���Z&���q����<3e�IS��5D��#ӋCt�b%ܹ�`�r��u z����U�&�-[6���n:����Qq��^��o�b�%�j?�kxS'ݻTc]�#M_9�tj'f��%��0��@��PA�ޕ��ۏ�JO�q�-_	f~v8��}��v�L���'w���2#ĝǮv��=`������@���+E�)-�+g0){���ܤ	�7�$Oݙ��
�I ���h[�͇#�B��6��K��Qb���,z%D�lR�VWV�o��N
�"�g�M���MXC���u_�Z���9&��$�x��6�����S%ŜF�#޿r�f�,�g�K]�PLՒ��%558��ïܧ�2��xf��iU�P����),�N��A���0���Éu�<��z�2�L���u����W�iJ	_Q��#�'�p) =Y	6'*�LŰJ]	�>�҈(Y���ض�	�|����� n�(��S�q� �`�{̵�R���f"s:��C:��1���W�aݛ���&x3@��+�yGT��1P}u���:0K��U��CUV��D���
�hɶ�Mr'q+M�S1<��a΅�$���|�rr����Ҵ�8ŧwyN+�p���/)�7u1��g���z{+Q���y�����sO��������qښ�Ų�`��ӊ�m]�Nni�5�M�"i�g��]��7[�#4EQ�m,��؜�~���0��
����F�A�O?:E�o�L��\��^�cZ/��L�?������(�|'hK�k�}/���ȕ&ʂX��*���x�B�����a,_z�� v���2�����V�|W���]Z���{.���n8�O31]<Q�@+H����
�� 
C+.y�#Ŗ�`,@F���0����X,� P81��j�#d��%>$��"�hB���:;��,�L-�!���`��@"ME;<bu4[���8�<Y:��jMi��uO�dt�u1w+�Q�?,��h��hI�f���!\�Dh�#���(���=�:3{H�.[nLXq�{ٵ*�<����S����^~�X�����٣ùB6��^��(|4��≤Yň�P��ߦIv��J}����ER�.E9p�������N{P����H�`]Q�,%7�-gk��S�ބ�S�1l��d�<~R�[ `�aE��e��<�}Y���p9bD|��B�R��J�6�M�m�G�e`"V�Y!1G}�T���p���WB����}�� ]�bdxӚaD8͒ڜ�m��q �,q�g��#01���mo��D�*t�ͭ��i�d77t���윰����;I�.=b����O�_�)����!�n�:t�BP��J&����A�/j��*�P�<�v
Gr��A�U�M�.[�d9!F����*��[B&�w��\:�U�q?��IK�qFI~���]z����V����CF���>:N�Da]-G�K�E��!�m�%� ?<J����t��)�[����*�j߰�I�$�����Mdy��"��
��J��t�<��H�5s5r���Q#W��q[bsI�����+ea���gB�*HZ�ܦ�II�[�)��}�j��%��X�o�Ǯj��?7��5H�;G7�(ۛ��f�e]cYMy<h�`�@\�R4��	@yP�TvhlI�W�n�U-�v�kA :������01�ު,4�e���n�G�#��8�#���'��Fg����EaΝV"A����i`��CΌ����"�������_0���+�\Я�FE{�e���٨�P�,h�Mr,m�%bQ�8��Ǻ~`m�S�"i��?d����9"�GA��Htj����������$�����?�8�߷�C�ci��N�b��B�"�aJ}o�𐋀�eFR7G��'��_���.��!a���eL����L����g[�w��p�7|�8�iy!)*9�d�=k"tܿz�I~���
qI�K\�$���y�_�o�f��7:_н�g���[���gM+&��_�#����ΙM��G�+)aU���%�p;'�2?������q�8��^"��xsgIb�����r7�w����9���:���I9"�]��:g�b_�QK� j*�n#��F�m���X�K�ʼ�7N/�;,�O�D�
����?��֦����Ŝ���mbUߊuhR��	��`#�&���4��Ǵ��XRA��/a�D���d:M��8�a�׉�9<λn�d���l�g�����uC-H���_hpq�cM��.f�5n8Rf6�?�$悋�a�[?�?K��\�l���,��C�*c�0
:-��5A���ܢ.ͩ]"e��}/���*C��깁�3���}�cht�c��������"�<���R�	�4K��&4�������+f�� LEC��4���5��Z6���VR�����?�p5�-^y<�&� pr���6�M�E�'vӳFu��c�i���o���=�����jXG���V�Ma	|�I���_0�
�jpr`�,G�[��8�ݿĎ�Q`�Q�[^4ͬղ�,��S,���tr�d9�)���蜙&k�v���g��(k�����f%t3d��S�y0&LwhbɦP��
0w$�z�܊#��-���8��9�FT�
�ك�k|���%�V����`�t�1��j�Ja���!�Ӯ���,�6���Ҳ��,�l��m)�+�yvn���tJ��pM���BVu���-���$VG��i��q�l� ����i���;�f$���h�9�_���ɡ}�9���?��"��=���o=��q�3�2/��f�H��������f��?TF'7 �%��$zJ�Z����j�}�8�Q�}WM�����s�	#�4 ٜ�A::W���w��h�u�,V�8	,P�\�S�V<X:���"�>8a@��Ţ/i�H�>swH�k���6�)��+mB^���e%DU-b4\-�Ȯ�!k�vE�D�zB���[=j8�V��j���y0�%7m�2d��=�����_���t'p^�5ޙA�����-l]�
�i�|�|��i��;��j�L�0U;�G��4�� ���ya��t�~�UW���u]�����Bs����b{<ϭ�Y�dW�J���+5d�[H���1�$��B#?�s�����'��n��X��6�`���ŢWP�)lE�uë����Fwh7X�M�R�O��zDx�:�Iw���sR�7�z�Z��	Z9�m��h~�Y����r��Kg;�;k'X�b����^�mCB+��[�oE�u�<�h�4�II<:�\�9h�F�A8��Mi������!�*�W������x~��I=����E��� ^r-#��%d�pEJ�� ^�A���[�����1n�E��P�YC��X&�<����[�oj��a�ִy��t��}B��<���ތ=�7uz����/�%+I������W�����l�"��rA��Д��Drm��Fr ���'Y�'��SJ=?�2c���3�[�t����r	vQx&(HI�%&�'6(%,�_( ðqtA��6K���g�����(4����j��J�ە�w�+V1�Y3�e�:�剪�%t�+ߚI��%{���Y��?�$=D{������]�L��"٣ך>�P�z���D7����
���Kњ#�YZ�'��WM��Mؼ �g�f��������\|ǥ:��*4�����0�f��#�)Gt3k�Hʛ�SF'4I��݋��0�m��r�8S�t�><� �j1�v�7y.���<b�Q\�4��"۩eT�|��^\�+Lˁ$�K�I�:�D�I�'�,� ��́8o�&@�K##�+������H(ra�>@�����f��Rj�>�4�V��P�	��ΆO�{��r�f��h�F��qңA�(���hf�v��w�I0H�5�"�����ޣ����0������k)���m��25a�k����$Tbo
3U� 1Ny3��	�����v����6od�$�,��i�"o�ᚄYT��r~����=��m�#���`eKP�a~�Os�葑dj=�Y�������D����]�Ȋ����N���E�B�ji:�X{*��&��481�6�n��-�5�c�w���]P�c<�<.2VMW&xLb�.E�=�_��w�q��4bM���ΞO�z�o�0
�4���քƮ�d�a���"���'�C�5�-��9d���Á�����!�6Vn�&m�6-)Ai�+�f��g��D�6%�����:��5�gJ',����4��QyJ!���m�AV��ܖT߱iֆc�xQ4�m7����.�`�	4����=6��������t!��]\Rϫ�G?�6_���إإ�J�5�#M�5|��"Wu/��O��6���!�/��v���V���D������@`��[r��uӺF�INN�?}����2�B��I��p��X��:���
혟����|U��:{2��ɂu����&Ş��p/P��~i�z�.F�8xZSȜ�b'm6��/Aڕ��Q?�M�=�Z�Γ̀�����vb�ǂj�(��̻�R�eY{욫Cps���� M'���8����o����cޒ��z<,���W4!|sx-Z2�3,�li�x����q���/?�c�W>rE0�I2���6w���;}w7�����x�y[�J����M�Rs%ۙ΢>;d�����a�a���A��}MpCX�o֪y���Gm�85�
![)�z(��у)FF�Ew(�r����Qx�����Y�j�N5-(Mv��1�0/�����*��$ݽ��Igf��X����cF�Z(U~��zӕk)�9�Laz��a�'����=`�k|;�&�=�uf6�Mı:=�s��79�i!
Ԛٽ�*�U�n�Zy�
0=i��䅩���.��3܏f�0�O�����d�!���%���Vޑ�s��_�$`Uo�=�5�÷F��c�� ������)��Ľ�\��8�h�]�w)�G�\�N#����G�P�V�X����%31�n-�umJ�ǆ@�]��Mq���H�����k�J��&��L�%C�	�}���q̊7�8u4zPW'��2V�{�r��������l���'��댲�z	��F��m}f���]51��-�\QIZ[7Y���zj4�����p������Rr+lK�V����W�h�G��~'��K�l�n�~�����*��G��&(c��&7l�v��5f-mo�����f{�n��m�	�r� W�55.!�O���aX�'��������p�ٹ�}'����l
�Y����:�mHL����A��3KƑ)�b��ԟG������QJ��V�X�?��][�z2�"�VU��vWot����=iJ>�IӔ*����H�N��EV����{k�%�ҭ��GWn*Q��A
Fpg�g?r�}|����G�2�&'ֹ�����+ x,�Ƀ�i}���Qn�������L����t�#}��Ц�̎��F���:ʦDq*��,��f~�\)��>Z�ˍ":3��nFn{�(b�=���<ى�'�5=�����.{�7-O�_���}(��l�u�6�D���ٺ���:��o�6��_jJ�r��ʳ����B�y���0���0%�6d�i*)������ ���G�bt��n]����c�����!�ә��Sg��(��%%����N��f䔹�-q㵣�+�0J��.
Y1N��p�ZI8Ƭ���r��s���a��c�-��{�;<}.5]c2}{�����Ow�����Z_�D<-;m^�DYom���&���@Kv��&�F���9�$�7f�,�3��.h�����kX�u�խ�L���4�z�^>��#�������xr�uIh��2�,b�B���<��g���R�^p���B��e=t&*\93�E�wKϷhhǛ�Kx�֨��{��`��/u*7���Ys�b�b_�BQyA�yڡ+n?�Ë9d��� �{�m�(�*u ����%wE�0���� O|#�2e����?'6\���K�
2ۓy= 색_~m��'�W4^U�r����4y@4֢���)%��t����a�*o�6D��V�s$�vI�Ve|*@oR8�1PZ���6�1Ci�C����ؙ��~I�ݱ����@_�ɷ��H��p���ߒ��x�ູ)>��~3<ku��َ���B��A�o1��/HG��w��;����0dL+�P/"�jS��g��>/0�*�����r��2ݔr��������\,���mv+��=(>Xh�}����ų��p�u�CH�w��/�-�<JT`�Fh�>��;s���<esX%��{of��@h��V(A�I���S,SN��:6uln�/'� �Cy)0��NɌ����[n���u��S�JX�	���Q�s`�ˤ��I0��B�Q��V�1븈�f�Eo����%�Y�imr�6S҅P�ץk�ӌ.�*w���u��7$�jP�B�kL�O��Ti1���uo��ʅR_c6���t�| ��s�;7�$|���KFm��ag�u��?֒������c�A�-��e��,o��؁IQUcp	�'���٤�X�����/ֿ �.L��j�'�%�y/����������m�j��j����,�u7�eQ"/���|��i*<8�����̈A�I���:�4$�E]���hT����9�+�3�_�y��NF�F�)�%.N^ �U�Xh-��465��øU���j�����P@���fs\-�[Gk�ݐ�i_��+=&�p��2���� �Ϲ��~�\�\%n���
�F���	�W�d�S� C�大� 8h�G�����Ю�H�� �32a�Yh]��M3k�G�i(��v�%���������(nD�Է��=>R�J�!������Xe�߻�y�j��ǡ��9���N�`p/�!2�
����I�.C����e�H��wWt��!��̒�н��n-Ǵ/�pS�
���YgUH������MS�l��yޑ��ʳb7g�!��b��U}����B@(��+oZ��'�ﻓl��Q��U`��  �k$�;B	������X���5�%V�>Ԕ�#�e�$�"�z�3�Rn��{ ��Ta�ܼ�59�%�6DՁz�ش��x1�]�6�Jy���%?���X� �[�٣5�
<��PB�3n!m�>�LL�X���K�W����]��E"_]��ܒ�)�Ȕ=���8P����q(�9�U�)m�?�h��	�*Er�r$�A�	 ��:cT�F�y"��H�1M���c�7ti�C���/�V�ǧ����z�5Ф)��	6�L6�������qP�G0&&�|�"�9r�P�������st���n@�p��
o��$��u����H����s�������*\��<���ѝ<)���iPLY:,a~7suH�-�e`>C��8��9x�5o�����,��KT�ؙ|�:O�;$AI��g_?�W|�6��g�7���7���q��/���a/8AdJ���aȴ�Γ'�q��t�n�1�#/+K֔X�/LBKEo=T��9�s�3�FR�oR��K؜3$vwQ�ř��J��3�pj�{�dPs���g�\��ޢ@�ܼ��>&V����N��)F��P�M������x�sl�&6�����#~s��ؚ�@ya�Y�0����1SF��j��T��~�O�=�GA����#�ܥ�[�sє�q��3����RWח(�[�]e����p�!_t"^S<��F����� W���z�
YU���Ǹ�^S�Xz��V��77w�_�;�ث{H#�WZW�/[H�;1�� �2o��҆]7g[ᢰ�ˏp1��ר��QT��P.'���>��`f����)weKag�I����?,�����F ��W�;���k������b���~��R�4Q.��wuYŵ?YtKK�lXZ�X���P��	+�$,p�sEH!\}J���F��a��6r�y a˞c��jA}1=9����t>L���h<8�7#	\J]=#m�RY��%9��Ĕ�±�^k��1j���bTE8�L�S���(z.�g>��0��r`�rgR$B�&��ݥ�G�ídt���`N2��,�w��[j����4��
��IXv���E�S[��$AJ 4�S1�\X�jDp��
���b-�LzKlb�����i��	dOڋ���{�T�7v�S�
[�e�+FF�Q�����F��)I�2 �X����vX��$贖������oǾ|n�%��z�.C�t��%�y�3T�������nؿ���l�"L���W�	*��Nf� �U��=/By!,��O�Լ@�2w2���-�;zH�c,�T �K'g����wK�}�&��A Hqi�MВ
]�泲�94�Kp��o���mc;��_�����7�S����3R�հz�y1M,t��	#U`�(Z��ۊ�"����D�xF���V�m����������C#��V+�>�4e�rv��Х�E��h/���н�>d���T�8���d����VI��|��b�Q�:B[T�8������u/�<$��T����貛酄�I� ����@���qI��&�G�*PM�.��ܝU����T���=y��ܼ^>01(A�6k��W �o�)��X�}}��%�5�,��!�K 	�eg>�H�N֋�F8e��#<~��Y�m��
د������1��;�?E���ƜQ4�#9`���;{^���ݛL����o	O��s2����	$��~Zf��C���i���M�*<��vz�B�o�Ih�g�*�V�r�#JA&z)��~H�M��ږR�u�219�\��nԣ�k�O�G�E�>+J?a�s�<��r�s&�]"Ǆ��m9� K2]��vc�Oa<���cN̓t̴��m�!�mv|�  ��3.K��	wvV��<ط�PP���.�-e'#'��9+�r�!�q�@�"���j�Aن��B�ؽ��dy��T\vgG����M��)n���e�GI��UN����W"��v�%�L[U��f�jc'���'zw��u�����N�mқg�̲*���/��2�Z�6i9^�#�@�.���:�\��������/�
�+dvmom���W��Cd�2|���ߕ�E	��!���}\s*�^/�a��Ճ�D��$���X�2���l%��Ȳj(�q��bsNǟ�d�yMz�M0�r�hsgzW6�~%'�^���b����7������;ҧ>��b&��H���g�c��B��ׯ�#����cD��?��B;3܉�wS���,�+#wb6lW���e���c ���s�``~y�%{��|�(@0����2�� ��:>��=h���]���v�=�E$u��Z��������Nt��D�������:�d�����T�>�g��_�h��r(fzR�lX���@�,^��f�}$�K顅|�� �E�CoK._ݴ-B�YT\��WI����h��Ɠ�/��a��TO�j_���:]{�4�:ҁ[{C������ON�.�\���\pq�4-��
u]gG��nS��'��3y����h�D��q֔E�SL&�t/���6O�����4���~}F�Ay�E�&��a�z���:�Xȩ:�yE��Δɺ�pՉ�	5Gq�_t6�AK1��o��_\��tص�^���)]�jW��6v�8x�j��uM�/�q2�.�|(�����Hÿh����6W�*�1��:�Zzp�J��"�4���:�:�kx)��� �L�Fx�L���(
^��Hj����.�
��%ݜg���'���;N�F��I"�}��k�K8[��L�	�V�ȣ�8�*���^��Z6��*�입g��Xc+SA�;��I�� Δ�i�%�b��-=�j�L.d8��# -��'��3)Zr�������}-^��q`j8!d���]���5Y��y֢2W�=��	0�C��%��U�ꇂ���v!ޱ$�Ba`�(�ǎ��5!1��p$������H=�-��m��oRk��]ۥ����ݎaID8r?sxs���9+4S>��d��G�a\�l
�Ƙ����X�rFj2�����8vx=��̍(��L`J�G�����M�.�п?,5���g�NF�f�om����x=��ʎtQ�~�[/B@G�@y*[;+�S���Ix�%����m��m�����ċ��nO7��uk���#�4w�D�y��9Ŋ��b��'�� ��S���U<���d(U��Ha.
8&���\��,p��;N���4���*�u�p/���Oh-57� /hR���N+Y1�nZ�`���Zꨇ��Sq��ݤ�Dz;Z����j��j��8��P�-~p���pW�`�L߻u�|�:6D�GvI�K_�}C��
��9�Das���'ch�3?Of�{1P��N�4���,���R�^�4Eg��֭K�'�X����R�s$�;$z?��nD�>�U����ń��;Ǚ�c�: Ñ_58i��@k����")���@U�W���:�f��'�k��)ګk�����17h���x�i�VS�x��¡��.�}d1�X|2R-�WQS_�������cR�b���m�,���� �XB).{EF��x��^~�ߟ� �Jin�6��gUjJ�cgs�]{��ڠ��0����<\>�*�PIlH�?���{+����Ǌ�� 7ݱ�Q�ѷ�_Ș�S��K��fe�4z��gD7kw�����J�S��q���ި�Q�q�J�a�H�T7��:��R>@��'A�QCƟCJ�+�pq�/s��E�m��>�y!�+��P�za0�K��V�z6?�+�q��)h�s�7�ᨊ�T�iŶ�K�M콳�:� �o�1Hej�&킳�G�z�����Dxr�����uI<��.���u~7�:H��5\�X�eQzrD�``���P�q�X2(�xJ����ƃ�)G�P�>pĺ�d��y�?\�u�3��"��<l�fX��nk�8�ZY�b��#���vPΛo���ұ�9�y��RY&5f�.��V�x4*����9�l$n&eӃ��C-�`�3�;�!�'�A}V�qAAz�� �˖uN6�s{�	�8@�&��5���q)��G��4��]���v��wa�ʏv�1�����G�����k��Í��� Y���	'jB3��>�������؃i�5�|�h�����x�
Xa΀�n�� �'3��x+�sMREg���kz-�����Ϋ�n����������E�NQ՜�_�^��#o�U����@+�GȊ�8�f3P�U]:�ׄ����]�G�g���x�s*d�	f�gF_�ګ���Jp�D�Q�hjʾ��5��6��v�WD��U1 9�<�Z���$	t7[�נ0�LY��C1҆�ls�-�"�Z;�NC]X�d"����$��wx��*ې�����tҳ�5�-*.�S�<�w4��J��g?AlՖc���(��0g���g(26���g[�Egu�0|_c]�d7�;~�K�9;��@h#S�����H6"g-�;WS������`eR�W����V��@N�����r���̥
}x���ۥ�P�`\ٚ�[k� �]ϩ0����:�M�#Xy���4�W�ܷ^�
Y�Lt
Ǿޠ6�榌��xW,�>��m�C��Ņ�ĘX?z$\��^�v#���^Pp�/�.+�+sH�d��(����I�|��tx�ۏ����p�\��>��ͤ��;7Oi�VT���7�q��bo��zx3dukS�e�d���f�<�p�ܡ�~���o�(�8���@%��.��u�$�u�vB�Z�CQ�<��+�H�j{��@q�C莫׿)^X��M�
��}������NF:����0w��"�y�D��Z��)8R���#�by>�-q��	����u��i�xߓ7&J�2���E��s�sw��b�V>�eTd��9yާ�Eum��� �h�^|��{�QX4O.����`��{z��q�5#*a�2&�t�T�o�B�u>o�y����'�
�e���m>�=����֨	��վ4���\�]4���j�:�I$�:�:� �#�Ԥ)�W�T��MR�w�T�B���+��k�W9���m��]��y9�x�$�I�T���HU\�V�E���т'щ�6+_��2u�7"�Z췈���_���*'l�q�;3P���k�uM��[Nk�7;tmEJ\XӹR���Hz�0�>P{E&�vV�>���32j
�D��wI\M�5�j��o��z���'�t�8�(P�;�F�4��@�2�C,
��/68�H�,�%`��c),n�`��B�S���Y�B��ϼ��Xr
ĉ�P�BI�j��&*X��n�wN������V	�����(�w�U/��w��ϯ@L�6�/?b ���$�XT�u)�@�ވ{3N8�ϋ��!V��6Ѩ�k��0��EB�DBO�1Ȗ��:cM��4�X�Z��~�s�N'��C�%u(!��;Ӯs�ӔH�?�߻�ne�v��%ʪ�(4�������>������]C�����
L�ܹ���f�}�h���;� �W�چ�m�`9�_��(���'R� [z���+�ilY��>�x0�����]��CC3�[���6�*�l�wO�t��HK�n�ǯ4VX̺��7
��,�����}���1���-$G#�O��ӈ�Z��қ��q��Z��Y�D`�]5����d���Aͪ��H��yU��.��L�&WY11�sz�_2��-�Ab�4�'f��Do<���oM9�Ϫ7x��.uv�W᠅�"h�4� џ���F�)2�.f�vyCh
���-n��B�I�1��$t�״-��M�Kbj�N���k<�Ւ����;Ag�IJ�j���j�s� B�.W�s0k�zJ�ɕ�Ѿ"�rͣ�Wz�e�����A	�����4��6�g N�g>���)l�&,��j�<�lZ掴���E�R��g���Y��>���P<���3Ƒ1b��،ޝ2���3�d�Nh������4cҨ�˰p��]Q��M�_��G�\�4H`
��7�	�z�nA�#��cB��6q)�}m�������q?�,��@�
?k���_�X� ����2� }(+�*oK3��C�}��~1:�4j�m5
J��s�q�p}��M���d�$)^jǐM��.��}�������UZ!Ť��m	L��wڋQi�j��9E��-j�N�,4Rn�u'�l�X��!JS�ܵ#L0��]��pü�������U��ʲvgZnH���V�x�������բjȢ�b0(v��.�����,��J�h(��j;T�M�~���P-&�:�ğD0�z �����ێ	����c��'�գR#��ɵ��o�(�t�S���������F�`�<�x�΁���0����O�pS1v� �C$�'Z�0�I�.0/AN���߶�_1����ٜ�;Cs�mV�k�f��KQMD&�gzW�oH6Ї�=�0���7S0��?���B�F�L�g�^Z�$�`*�붔�.�G�����/��10YFk�뚢@X�ա'Y�2O��ΡF%�x����n׭gŤĚ'�x#��ynY�Koop8{}��9=5�����qV�<A�р.c]L�l��FfQ?s�MQ���������踤|&������T�άG�#9��`�t��?�ۜ��0ޠ .XkC�eh����	������y��x�����=��X��ڨB��d��-���"��q	��~���U����h:��2�Fg1/�ʑ�{�r���d�_�
�S��?��3y�_ܫ}�hೡ� ��P7�➍��wwm���c���~��"�����~l���- ;8j,ء��z`ԛ��P|���J)u�;�T������a���5�N���|$�|�_�'@�ԨA�gB4�3E��̓p��E&�X'J�r�i� "��6����5����G�Y��'fn�x,<�L�U5VY�J45y� �'�Vj�#)����̿(�P�*��AG� Q�O��
ˏa$�N¤X�,�������ݶt��k�Um\��ԟ�>��x(^��~�kv�0�2`��i'�~̡��{���1�Ƚ#��_�p}^B�[vZ*�F���E���^�;&�: -W�VO�b�t���� �C�Q�S��G>̝1utt�o�3���\��<�|�(%Z1�v���4wE=�wצS����FV��iWO<m����٧�Fx=�~�p�sy�b�o�@ԋl��F��z'��/��1�b�a�cx?��Ť0/��%��u��y!A劝i�=�L���B/��WQ3�%� ��`����PO	��#�4E�� ���������qz���"�n��L�}�F@��$�6!_o�9gW�����m�x#�%GҪ��3�qvx	h�a7���GS&�,�B�I�X#h(�w��l���NXy��צ6�@ö�e-�{�Fq�*P�`~��Y6���­�cʌ]�W9/���$
b1�ĩM���?�"џ��Yy������Y�w�")��'b���T�wOuѵ�ېrn�{�k��:�ǫ�Kn��~e��x�T�}���M�v#��K)	>1�^:F�ʋ��$�ݔR><,�{�4����tdzi��xY�M:P��2�L���3��3�S����eR��wl�џ�G�#�b�t�Y$�[s��Z�Ǽ�y���������7p}�� /���O��%�n�������$\b�9�R�+��Q``W���{|�\�N�v���!�pm�����(% 1�+3���mԒ��y�$=�;�3�N��=�����E{]N� �9a�.��������k��RͩQ[�U��*�.8&y����q���c�j%�/�(^�8�?92m�s�M��V���$����p��g/�w�T�!���6��؇�����m�B�&��֍��rw� ��>��:�MStP�-=A��Vy������s�0^�x�#�s��pK\����E1P��l�Fs��D�-���8u�*�^�y����\N_O�(��c`�g��h����V��:�A�<�KMȪ®R��"�����07�ڎ�0���(h��1��ܢ�vW|�LU��Ϲ�g5Sn��5�arjÐc�1
Zf����D�\`f�D��j�K�&�=�<qn�,]�G��=G*|�Ш|��x�O7+4(���G�A�'�~��xA�į�����n)�̳WV��:�`��̊(l?����Qߍ�]^f���Џ ��\�F�݂�n���ӚGT<��
�e�㎏��Kۄ-��9R����^�?��Yy!��������6r��sz�r� ���$���b�^~�H���9G�GAt�����-��O��:Qͼ�)����{:��"m��9}S����yE�W9"�k�����֩�D~�]?�1]Zړ���䣑�:򫥊�Cѣ��i��W��j���E� =�D�����.���BQ�c\�4
�+�2���C��D�kќc8ˎ�+�̏S�a����c̶���Կ��VO���/�Z�Q4��B�C�4�=��Ҳc�~Kc;��W�� ���Q�4!�;�� 2���K��E�+akK��9���V^��������FS03*��s1�9��ݻ[|�!�>�27��d4�� �v�n�*�x�CAï�K�g��^�߃�3=qc�fĕ����Xf�U����mS�PTf
��V���v�֏�I�7�s�8?lGͤ՝��@�,ܸA�\���ˍx<-gwk�_�u����JXđ��Y"��D/_ޚ�ݧ��T��-�U:��̷����X���۽����8�z��h`:�����(���jk���W��y�/�٘�ji=��M�bH�K�#�TV}�yje;�u ��{����6���ư�|��I�v��ֆng\�E	�H*T<��OD��R��{�lv8�p4gX3�0hf6V��7�q�T�s�K&!�j��zg�ˢ�?HW���#�ڶ����+#��b�[��-����P�kv9���������7��������fl�p�Q遯�y�dMj�E1V�RY��#�����7 �Jg06.����|�P�=Ʌ[�����*��wu�<�p��o�"�3�G�[��2k%��41
�9xl,k��h�k�z�<��fٌ�xI��x#*��f�g]�'���U���!s��Gx�lJ�Ĝ� ��F@�5�ul�� sco&n�d�C���Ң�	8���l�n>K;����2�[�*�� ��h�ɪ����h�(�0��"AQ2��c/xC��F��i���6�]3��L[,�-"S��v�' �\��X;�����rļ2�`�8Rڠz��8=Js1S�b��%���,RF�X����NF��
�o}�F φ�[C���.8�5Ut@$OQ㈻������y��t�;	���5�M�͒���4��(Y��(����2�e v�`���-�5��r���	~�Uw�P��H驧}\IΊ�e�u��98��Y#��ר�c�Lab2ɡr#P>��~�+c!d7(}�?n�{����U�.��LR?�$���B�6n5oڐ��=����N�Ϊ(�=�$�qg�nHY�]��UV�t�O�*�������M6.([%�ؿ�ϱ1
)���`�6�+"�]A���_�.��R2�����\5v����^��C3��ء_j8�[��$��pc,q�����E6�|j���^��T��G��� ��At� O��N��J���Iltx¶]�*�wɡ�ډ.ƓEg#����)�d2�Ё�� _����2���O^��(E%�>K�,;c���
�J6
�,u�m����;��J����?-��B�C��<1�Z=�-�"_�N������D������'�7w��RO�22���|),)D����͏ ���|�-娑�6�!/�]�ˀs�c�kGW&i�a���Zx������7���%DMI!��2��/�9���!��i��MUo6̴W,��r��D�_RY�-HtF`Ѥ#2�$��$9�����5�ߞ�t����o
�%�(Qo]J&?�q�f"W���(tUtT�L����:��lx>�$��{���K��}��˧��`Κn�1-�w�'�c�~�e�y��r^�?+�)Z�~w>��z��WU�B٦ i�m��U���:bJ�bE�
m�qR����P���M�2�?.�`[Y��Xg���JN���y���8`�`]f,L��#n�t�_i�5�0���O�G0c�Ԅ����id���Ȯ��3���#/�w Gj�N�F^�+�����N�ñ���.��V�-B4{���FuW�^`O5VFѬ������,�n\a#|�z@l:����a9��5z���P�W�E�=�^@!�**1�a[��z-������O�lw�M��3Ox$*�����*��[�MدD�M�By	�KB�Ŵ�+�������\�NeW߳��&�ԍ�z�+�;܏�fs4JPFʴ���/��/M#dx{��\٧���~hN�USF�a�ޒ 3۝
8�θ��J�u.����VU�)�+%�e���M�a���=У�\��g�{��Ĭ�.�����l���p�e���4.�}���k���*�����@�,�3%��Óf���[�������_�*���Y|�{��-X 6��DU�)F~�;�U�y,/�9.L(o�}>�{�Z�(t�9f���0�����T!U	��==���\�߶-�ei���<����#���.0V����j����[��w
̦��gm��l@��}ƕ4[�B������o�|���gXT.3�<��Xp�7�a��x�c#n���-�����B)%��N�f���3�jf&V��v��{��p_>A㎝�t�I���Wc:�u79�[��d�F�t���]��᥿w@2j������%�f��{+���Q��g=A���n��Y���f'�Rbǩ�N�mT�{�V��� 9H兼�6�3 �Гd��C���h.��]t���Dl�,���iEB=�7"��n)�o'�P`��p1H-+�cW-Ⱦ' `��.>�>�$�2Y+�����}x��f�F�ޒ4�įz7o�_17���]p>�7�wҶqp��S=L�q ������e=��6&el7\+�1��Ð�p*���؉a���>�1�n�R�ح�����1K���ɨ���"kJ1���t~���>��&[ d���|��6��ie�����,�Y	|�%���n5�i�Ϸ��*+��W	4��"a�p�����-���5.���M�0D�on��Ì�X��ǝI����'j5��� �\�D�13B�;��xbǙ�`�Ƙ�^�)��R��<�~=�!��� ��2l�Z�n���u�u��j�yFS�,AD��>X�"�������әP1���ێT������������{L�����;`^�����]/a�!G��d�1�bM �����j�Skԇ��( u�����C�и̳�+Xb���&4ەj�<����Y�^�G�}*��ɦ:Q9TSngQ�I4�{�lj���RT�rhDSd��Ua;���`��F�q6<.i�0/13�������ېT�Ϸ��yr�y���k��a*��J��,~��p��˟��;-�\V8�s&����$ C��Wv�'�d���F.-���p�'���s�Ԣ[�����2Ĩ tl�	�5���t��o9!�3���Dqw���ũK#t�5;��%����8�6�Z�����{�pYg��~!��J��x���Q��+Zm�<M��+�WzV�I�߯����� rlޒ}x	<)W@��BHSq���)�R�~R�x�sm� �MD�����<Z����u�d`�M�e}��y�f��e�T~��������Ģ�ӣ����]K�k 3c<z	�CA�뚴rX��u@T}ܞ(�U���C"؂�@a�cĨ�-vy&"լBa���?��P݋Ie�6�/��1��w�����vK4�=z�f�zb�s�� �|.�@
Ѩf��]����K4�{�߾�B���ڒ��t$��A���7q���A���Ī��o�=��2h���!��Ng�,��|p_H
��
g�6�5����O�9���?��7��!�-�.̪��b���טƄN-��hiYt�,��B3�B�C��^\E૝,�Ю>ݯ���4;d��rC\�b�&K�'�xQV�L>w$J$wE��Խu/�$�����!��ݟ�N��zY��p|�zπ�v�A?�ުX�0=sӅ0�;A<K�?}řnn�<0,����It�����m3�,���J�	��t�#�V|ҴQŇѤFQ9�ɝ�Н����F���
� 	-�@�;Ly�M$��	o	lUߞ���ԅs��XK�<�=�ͺ�A37}�o��3�o��H�!��i�.�GxAω� WH�`"<8�ҟݺ�t��D��Kpuk��갱�-���kT�K��?ءj��0\���i�=��7�-�����)�g}u��6��a���cd����!�K���#Zv��D������Taïs�sMX���<|�]/�k.,�v�B�b�U4�Lj���ˢ��./�l=�/}���SY��������!բ��e����8�r4b�����2�"j�l�����L��8"�O}F�\��X1��;N�%P?|���5DN!����a��Ĝ�㱅a�{�_�s4M�ݳy�K�:�Ag�����<�7%��d�f�����;��B�}���������๗o7 �钗 �EE�h��u3ؽ���<W�r�FV�i9����ǂ�E�~��0��_���Oݗ�)������c�e��
üS��ц�S�h<���hc�7�|�[��TXpC�Ft�;������(y��,��@�$�ؽ��Pb8�`�#|�7��<��6[:r�Q���t�������M��l�DO�s&��7z�V�q5�c�R�􁴧��H��VH̵��op ��@�_)-�꾚�X�0f�"{
a�|Ê
\Md��O�4qӶez�����$�$�Y�}4{}`��\�"q�R����hяi���t�wP�/]����Z��y��`��fXSq��`��#�"V��T2G(x(��i�Cf}�0kh�g�C)�Q���O����p緼�3v6�>�@���9�=>#����f�Er��w��+<����,�/+��z�;�{}�%��@/�D���ͫ;�6J���P&��ά'E���<��o�g�3�2�{@���>qeA�D�v_XP�%Ȥ���j�Z�ϴ�s�V.��a,��?NR;��(H�Ԝ�Rs��բ��Ñ��ќn��[���n�����R�vGLV�)������jG�	@ȿ�.�`'�s�-�k��5����|�&���w�f�w�g�5o�Ӂ.����'a��ٯ�K�I�.�����X�tY�L�L����t�l0u�m��M�NHf��'P�D�M�K+w�Յ��)D�6�4��fkGG� #$����xցB�uQ�X�JQ[ߥ�bЅ����-�!��y!��}�J�����Ǔ�	���D�p��q�E�}�c�9�޺�E'��T��%f������9Z&��D,}�I�c�̝}�]��9�����@t�&�����L��N�Fɣ���b�����������q�68�V���n�UE�>kgwW/"2�M���}D%Y����Z��TA�6����}�{4D�����<U�GM�i�?]E�����t*���_��g������^ t="��Y��P��9O�kS/"=��yY��S]I����L�4QT�0��;\�dYnp��AX�W�,k���lV���S#ϫ��izc���{ �� w�K�������3`���ֳ�����ex1��I9MT��g��rP�[�A�i�u5�7'�_TrLݭ��K��+|oNE��P6#�)E����|��9��.���E˳�"��T%@��T��U=�!��~�V>�k��n�L{� ��!�?�0����g(Oߪ!XD;e���v8�o��3MP�"��R+�^}P6U��r>��D��h��������mF��`��1��FD������cf���m�R�]MH���L(�~�x$ 1���0����DiF��ip�]⁃Sd��H�� �#�;�1J�!�ͅ������R �x�u"&�Я(ǘQ������,G� 1�bG�ɼ\�s�+�`�X��gRB���җv�Y�؅	���b�/����qJW?��I���
�
�k�,��~"gn�"=�a�]/��'=l�x����le�P_��	Q��̄<�f!�З�QW�+,�b����0S�.�4T`���e8Ӎ�/�R}������C>��pA)�OG�����	��Y��W�n�V�nӟ�^ΌL)t��:���\n2�w5 :⡖����m�-.f�<*��ҁ��V�a�B��i���b{ޔ���2/���	�°G�����?W�����$��u��@�cj;@\++��K����V�eM`o7oH,?Ix�a$��q�����SQ�:�t.453_i�����lcf7$����H��y��O����Q��k!7������CK�k�%��"i�x� `�>�Y�'���;�D���D����>��I�$���y�ǩ�{��c�����=r��o�Z��o��.�4�킝𳶾���T�肭����o�պPn�)M���I�p���'0=.�i~/1G�N���O*���nǩ�sɪve�d�1�r �P���i"�f��ϩnwi��wh����jҊ�n��a0�n;����c��b�Yъ�[h��J@o\��]Z"x�׫+db�,膿U����'՛��
��R�=�;bn�+�z� �bc�BtTYҭ�d|�h�ۻ��SH»���o'FOF�<7~85��l��q����³.	�/|n�q��W0O�6r�z�츚޴p���yo��g��Q�H~hp���[�I�<�a�L�adl�M,�{ȴ���� �׀,�⠻d��[���*���zDi�~z�
	L'x(��"���MN��*����嵝����c�"��Hp?j�f��ljb�͒ڽNϜ�ӂ�/�-��pI�Du0(K�R��o��yn\Y���X D��Ҫ׺����w'��I�Z�-Oekse[I����>�W�0D����:,��~~���>3{I�"+�Y[S>�9�}�D	&�c=��.��s����d�����.4Js���bp��w�hs��pt��:��o�<���o�/�l���������7��P=�@X��ZY��?y=�l�@��R8]����]�eM�n×����� �pi�����K
\�b"�����]�R��$����Ej�Y�L?��s�ܤ;���D�b�0p9���`ևݯJ1�~���a��{��L��Ŏ�	t'T�a�߰1�*#�I;� ��F���c��o@���;���8��3[��>��;3s�\��:?C�Xu��@�.�db%3"�@�p@�S��w���mV#/��iP%��{�a��"$�uTQu1\��Ot�p��f$�ܫ�0O�~z0�_�m�Ҡ�+��T�
������q}b�H	����?ez��h�$ev��fc�k$�q#�
��@��.�"l��G�4�.��c�:���t�5���+Q�Qt[�m������A��ڀ���5u)p/�M�	�˫�G��t%8 ����z�=)4B�����!k~�����32��=�5J+��^�� �B�%yt�ɟ��!���TH�z������.�o�A���M�H��V��.�N��=Ū��PSGn�@�x$��W��As:�C��D�k�	���7~�J��0sY.���a����7H�����W�^��==�xo�M�㑢�2-Z�Z����F�Aly����;��An52h/߮���1��֡�Z�,\S�� ����/���z����a=^ˑ������򒺏��S"��C����da������������mB�:[������mQ�N���\�Xw�e���ۀ5���֟Ok-_�������G�j�iE$��ϷM*������4�����7!�bq#��|$٦�[�-�.xt��[/��V;Q���͠��g�^���R�L�~���(p�|�i��q<��"����n�3~���4xS��ޖ�&k��0Î��ZLacϺ��TX�\ �l"M�ݚ�u2���#rt�ʬa���0A��e.P6��YIs�0��N�"��)���#q�����ӼO�<�	�����](�#����������OsS�^��%t�ȷ����:L��W��.�y`G̦��a6U�����-��M��{iP=�j�{&�y�S<ꇑ�x�۾��Ք���k���B���,3���B�����GoC�&B9ad�f�fU����Gm�Yͥ��[J�Mަۥ?�D�!�筇v��7+}2i���̍�@��_�T��>�k�C:Y��mw� ʄ�Eg��P@��Iu����<��f�M�C��c��ޓ�f������z˷H�w<��e����cp+�^޺�?R�YV�s�W���>3�}d_(��ڐ��0���*�ےO)��[h.ˈTaǘ��.w���I��)�9\L��,�5[?x�p��M�d��Y��%���6�O��^��-��͐�h-�"o�@O�Ƒ6+}�(������ol�z��Cљ��y
z|񦲚�ќ�l�GR(�F&6L�К�xƘ ���D�̕f=n�O�O���ߵN�Fg��3����p��괙l,���鮿�}�����i��M]�$>T�Y��H�|(����b�u��1�U��:j6�@�E",��~���\'z&�,���dS�z����j���7��Ї��M{���f3L`~Wr΢���0�H�Y��#9��ۻZ�<��%�1��� ,�]����{����{Ys��WR���2�}{�1�	��u��*Q� �k�&��+͕��/:��awd�a*�\	�g�+�K�N��/���F�����h�j-�����=�Xˣk�;��ڦ!�9��,�A4{����˒�B�l%ZL�e��ظuV+����F�[��������v��cnit{q��;G (��8O��r������ .��c���w����0�V�H)j:���6l!#Ir��*�E�H��#�3�z�}�V�H\�N�+Ne��p	���2-0�$8��G#�3�?$��/	K�w3����S��c9���HH;A"O4'R[2P�X�Vo�j36P*������9'��<�R��.�)�Q0Ɖod��>�,ދ�L�PQt����=)EMiZ�>.c����4�����p�7������T�D��ʖ�,�D\�%�Z����r���"Y��?^���A3��������H�I�金1+��z��q�v�q�FҴ_TI����y{��L��v��R�,����=7 l�{���6Q;yJ%IRQ!���p�D0.�mmw��*����Ti���qt�\�/#L�K�UE�K:�����,<?���>8A�-P�UL���b���B��v��G��՗JzI�y �"!�r�<�����WW�w]�v&�8⋄\@�>��I4|.+3��U%�֥Gح_�3讓¤(9���n��H����c�Xb�	�U�2DR���.%�b9v3���|���2A�R'y�ɏ���^���P�Uq��RJ���e��q�SzL��,N�ȯ�p�����;�$j(`�,��D<44S��;+SŻC�D����?��@�F�k����\�p��>�V8Si"����"������b	� `�^2�lK2q/�Z�aJș,@��#A���%�����8���8��;��L�������c���Qe
D�Q����wQ8T #��[v�o�ԁkf(4��NZ⭔Ԫ��Ѣ�2��1K'�2~�귅�3X�����4Ih�.j�O��hL����Uۗ�:5p[�%�߰A�,�P��?i���?y�jG_�]�U�*�.p�F�u �1��D.$W����޴s���v�8{��,\���a;U�W�k�������2���Q���bk'���
����7p�{�9.9�l:_\�#�]�����|�M�:UZ{?M�P��]V�}���P�cZ����,�
�(��ހ�&=�o���Yj��Ʀ�%�+|�?�0)��#N�t����3��7/�-]{ǂ�?|�3�6y��C*to���]O��]y��� ��<`�d
�
%wQ.D��<�'�Ǉ˭��K
�b�ACJ	�V�����^�r���?m�HO�-����ȟ5�Ʈ��3�sd�fQP����������m�����B�������$7�l�#~��ŭ,#<�Q:X ?�z����.����yNa���m5U5_�A�l���+g���W�<P�J�QЌpu����E�d5�������ķ�g�ZY�CE�%hB�sXi��UA9�vmܴ�e�H7�I+�Y��$D�G7�
��I=�����~�;(0[`��������(O٬O���7�ì� w1{P*�X�-,��1���S���NE�Ȯ�rJOGG��,��q���Tg��G��Nt�iX��جS��/��2n�2����o��+���cF�(RwK��u�eJ���x��#Ot�t����|Ij�VàQ��S|��R-u�1�|��v�	�����B�`=��"�Y�<x�X�	��|[��aX�IN���B`;�����ȍ���v<�ۧ'<�ӛ��Ă\��k>���P�� E��Щ���y�S�s��r�� U�g��6����<s.��Ȫ<��:jmj��Bt1�������=
���ƥ�C�]BH~5�3���䅮藩�
��F���e{:D_����͉J��x^ul>g��{^+g.�r���'�YcB�S��N�r�hb �n�:�oi\s����y^u���zR;�[_�̌��G� �l�(R~fAt���҆�p�F%�
��;��^�� k��?)��:I��ZW��~��Ȅ�\�R���.R�l��KEp�}�����{�+�Ϗep
u��C?��9������]�O���܅׸Vh<�A�ת�|�٥e�W~���ހg���W���J�տ諈�g���F |]�z��<X�"$�����эl4��H�K���R�9ꫵ,�=?c��Z H�N���+p�a�~}��k�|r�AW���~�X>�aF�I�T�s��X���lű�4�{Q w|?���أ��%W��x>z��E;����r��C�t+�ID�t��'�69�ݔ��nlL���BSu&�"_����"�e;%�^�
���;n�����W9�=�/9�궩�nO����؛)z��B#��d{3�?t�AB����q;��7>��c�xW�GkD`e3�LBt�� s�Pg��+ ��1챾M�|=����Z��.��4WCR+[�3f_�� g+м��K���N:�F��2��X�4詘������9��n�����U4��'�i�L�����q}{�T����;M�"[O���7��U�A˿��T@�?-�g��ew�x�qQ���ҕ��C�o�~���"�[��
E#�$�7�u�z��pO6�2���yq~Z���\�Q�0���&I�vN�vz��`��~��v$y����k����|*j�� 24�s�V�ל�?3\���oXzߥ�s^�/��b���⃚���;h�����D�1�8���\xX��߿����F�n������v�9J&�Tw�B��Փ44p�E�/ؚ�+,T�K>fH!,ΞR�f ����H[m� �C���}���9�sf�hn�kS�9`�l�%��H��uY���s�@	'c���5�YL�R|�j~E�"mj��ma��n �vHS2�-�F�25�*Fr���E�o�7��t����{����`��EOê����UM��v�1�$\ά���D�Sᚪ������<�����]"�W��Y!} ���*��K�]��6��|ۆ#�E��\��x8ܕe�6i��`���CD-;�n8�ˣ�P��=���x�ek�ʎ̣��)��G�)�C�x�0m<߃�E�k�`$����v>�*�?Tԥς߻p�>ݔI�1lL�?�W����D�Lݓj'�"�O��ɲ�S�`��`�:�� �y3Ϙ��ۏ�ّ�8��(V��|���AlA�~��U��B��n'&e2��$�B(:�F�y9��{е��؝��8^��J�Y`����W�R�u8���zE�I��-t-�{��/�)�]�n��I}uD�n\k}��]�S�%��8c5V����ʔ�ۄ1�O�����n��|��DvE�4�P1��]�*ae��X1#��Y'Ko�G�5�s��3�OЪ��q�O�D�u�p����ؽ�����{��lg��!^�n&j�����/������,����Wf���l��;r���\�b%�	��yw{�F(g��=9��F��L
�QQ����M�O�\�#Q�r���*p��ډE*a,֩j�_C���"�U$QX��N����h�@���D睊x���=Ր����дV�*c�:��X�~�	YQ�^�ꄏ�4rY�H�dʖEg��8=��?JQ�!�;��T��y(Qe��ƸV<��q��|şXOG1^y�h�����3�+q��m�Z�f�9��EA2A^�fS�as�'���`�݆#��j2Ǭ½�����釔}��ԕ��c~����4���n�֍�-5�h-L�/C���F�+s�A�~�]��@"Q�	mu�E����	i���BJ�� �#p,ۭ9��|ଉ���#z|��Dr��6�ND[���W>�	����jZ�s̬�ȫ�B%�lW��c'�?�K�CC��i�]�"������N�� ��o$םWW�Yt��}vO�	��w�@
�g#��*���:��.��R��o�����a-2��l6�>_��0}�IΗ3OrR8�a����ۮǼ�\U+d��:�;M�Mg[��-A]b�3�M	�_�Zii�c�n��(7�^O�@����l���-ët�A�jD(}��L�BgWe��~ 7�}5���|�!!��w&�ڴ%3N]T-�ƶ���J��� ��:@eP�K��L�|�%�yj�J��$y=/^�!Ic�������T��P��AR��R�RϮ��P}� ��c!w����l$��)EJ�V�-c㨜t��*p=g6�������>���6�Y��uO��WW���s��	1R� Θ��0B�4p�/����˧�Ѩ6���@�Y���=�RB�Z��~qipF�	JNN���CźG�T�"�P_�Y�/�@������L�j[�D���M�~c�+�^y�v���j
[�+F���C�2N޸���N�LװOj=����O�qT�=�Od-a���sLR�~�\d]?`���N�va��'C�Hl?����v�zݣsa|o^)������$ބ[f��K���S"\�B?��C�e~�o�Nu���(8�%ީ7i�n��kIZ��߿�o�n��&���cg=,m�z���r��NW3�I	�:L_�)Լb3���]���~��	13���7V���ɬ�q����fY���9z0^y�Ē05"? ��Y�<��b-��\խxS���^��u��lx���oR���Hr����s��"�҈.O$�D�n���Lnp����&��g� sVz�wBU�<�3W�*�����a��A����O��dW;���v�;�"�75}�%a"�vO�
�&u'�,A��)ڻ<����D����Lmc��]���kL�JI�2�P�zA~��qi�����v�\W�V���B��%��c\?����	9��Q�RZ�e�5�1/^(@��3i��)�-kӠ���߀�	c�A�?�l%��v!5#Q�����	Lb�'[vQ���C���]��9	�Y�r�T�W��堛���G!x'��%�2�v!����xK� ͬ�#����'Xܚw�V \��	A4�FƘ)�9^�1���J�����&�>O�<u��U1"䆚G-�K�h���~S5q���2 s������?Ldg5u�Ss4i8�2�Mڣ�k��w���'�g�F}$ZX#��^��AճlY�wߦΏ"�%K�b�A�J�A����D�s�EYiQ�����T�W3���\*�~�p�6�#��"�v�����U��QЀP��d�'���w�u?
�u�~�}�����DU�8��\S!�,z������:M��<��@o�3��Os
���~Eה`�f��X��{���� ���9�H���GD&pK����@�Y洝CYZ�O���M`��s�LI�3ޱY�c#H\��&���f��"���U�26"y��Yl���?�ޅQZ�v�9]������9���t�(xm���w��j�U��aUWk]�ku��߭a?���Z��_���A�\𧋦�ԡ�UR%"%]}��5��	�X���� ���>�AK1�ޒ�cv�nA�<��l�����R���o粆?JFêwR��=��ΊV��n�?Ԯ�����A���~�ٮC��m�ٯ-.W�[�E�ݓ����.q����*m}!!��;(�	��:��~젶q�������h(��CJ$�򶺅� _�L}QJ� b4�gG��N�Fԧ�i�\��}�&֢� ��BJ����\��,�$*D��
���w%^*��Uhx����2�=&�s��)!&�o��O� �]?g����d��4��x�lh�ϡ
�����~m�O驦6�6\���f���G� �e�{���ؾm!��W���Ύ���l^~"�[��?�ᓬ3��A�2��'#�F���tpׯU_t�2�Q�i�h?��F�(3�m�uHC�*�%B�NrA�'}�=|��'�,\����	b+�r,΢~�SP��'��^�9��j��Ԝ��t2�D��JnL�p�Tuiu�z���j�2p�a̓Y07	s��DzK��m'{F��2�fꚵɦ�p?Eе��+���Q|ȋ�*N6�����7�rx{���'�?�p���&?���S <�X|�wGZ�/.�zB�Հ=Q�dod�r1C��qq�1-��Ww���J���X�fu�JkՁ�I��J�_3}^������/���Hm�g'�7��E@��M��l>:#�"
�N�Q8���H���V���Fё5��8Ҝ�4�k��s�aS�U��T�4Ϗ[3��wo(N�Z$�Lu��/6���5�*2���&u�X�x5�w�w�<M~���<�1��Co�Y��L7��e�%�*��;�❭x �e8�?��y�������<(�$�˧�
�p�P���G.��"}l���?��p��uK��Q�d6�Z�
�;Ц�Gm:1`��z4 ����L��R�7���{7���	���%��c�_�?��a�,_s���gy����$Ő��C���>zI&Z�F����o�a��*{e�\��7���WE��ٟ;
�Z4M��.�_��z�r��|8��@̐Mh�]�dg or0�O�O�J��~��� ��� O�,���M�Y�׀x��<t���?��v�BރF������j��߹|�1G���Ǣ'}KsX���*~��q�� c�)QyD%��������<wYO]tgx�lS.}o-��L 	�K�7��t ev�^H�Ot\��pt�GJJ�>J_��~�Sch�gQ�����=#!$٫�Ra��Яa���<��N��G��tR���I�6�3!�$y�d�I����j5����r(z���x
U/'m�s�A�;4VP�"D�Y�����/�wλr�t<�������2(������a��)��Ӓ$����g����.^_��*!� GI���5;�]Լo�(-g�M2-+0-Tu�܃^�*�'�G�Օ����Q�fcP����M#��=���p����Ŵ�y�D@�P�����~s(>3��R)�[���l�]]~�s1e��|y��^�1��߾��Ȇ�jBc��Ƶ��gLrrV�uB�xo�+�Fb�J�ϼ5���a�E;� �h\�ɗjvH�gǓ���Oл����u(OL��^Z�Yaa��Jx�=�|��N�fMǅ:��T	��HFU�m(�} ��;����0K�sƫ�_��(	����biх��.+m]�M>�K�'�$�>����#����j�<��.~Z��1�Tc`�y �Duw���g��w���9�0��f6*��	���HK���%���	F�a������!3��i��y{'����_���I��G׾����:�l��Wƃ5��tOOM��_���i��ze	�TW�A}Y�,�T�l,PbAV:���VE#A |Z_6ͫ�m���c���1� f���E����g���u�����?��q���B�9��oǲ�A�0�[��� ���M���\�*5�-h~��C�[��
�^l���.k�<#~��X���E�u�g�z�sѷ(���6��o���Mm�F�đ� �,z�(%BĊhE	QO^�9ꜙ���u(��<���+�Jp�rλ!�q3wa<����{�(��p���{��>.f�����yl��h���� H#��q�K�҇�eV���������DʛI���T(D5��Ќ�*�l@v�I���qFUO��?wc�2"uwғEt�8�Xhǭ�],Z��]���9�C�}A\����߶N��%v�|i(�br�@�(�A�媢��S�q��E�d�G}���O1�/�Y�{�U�mf�_Pb����߆Hh}X���F����?ޡ.7ñ�g�+�{�yͷM�oJ�����#��ˊ���գ�$O�=��9OP���U��b�v�M^�ۓBV�(�8ǲ�nd�,܅��\�39VS�p�Բk#�x�5���U�]�w8�p�2�'ӛGvׄ���<^Р\�59���<���q��?w"��;�� ����Y}�h��s�?S��� ��*H�}��@��7���]Vw�t��)��׼jJc"!|�)���n�pN�3
;ֆ�|S���/¦{s�mf �2���+h u���A
o7-�]Aq����sEම�#����a�mfN������8�*#��/����� �Y�,�k�gs�&qA��s�F����Y�uAB}��������'��S�%F"��cp��j0��O6VQW��`@�yXs�0�����s	��,9�{�IQ�~l�z>����M�K��@O��ʄ$� ��1��H����~9mx&�P�ilУ��]fPʦ���C�j�3P���-B�M4�>�^��8G��_L�'+�0�>s���Z�8�޼�M�N+l���=k�Wg9��i�
{�����'eh�D����t��[҆z����}u���Y<��ݝ��!s<*�)+�6���q�傗8N���WWH��j�
�E����i*{��Ӟ{�?����A����N�wR��?�d��X�y5F���,�Vps�;a����Q���˟�,����jf	c����hw�^����.sA��}�u0�Ne����J�u@Pr�»����q5����BCv�)?�Le�E��Mh����%hc�{�&o�l�L��(I��y<����G'+CW�ּ������س��u���Zp��.>iC���&�a���Zl4���/Z���b��EC����\�@�f�Դ"�:eR�*�(߼8nO/��;����P<�kUs����j,��
�;(��ޛċ���f����K�
���S,��>�n��A�����9(Ԩ^'ޓ��S>���JD����`�5DWk7󫽇��>�A��Q5�C�>��6��C�01Z��`�]?Fe�B�fF�EBQņ�=�ǐ�u���V�	�F�[	C��. ǉqos��Sl� ���B�*9Up`9�1_�&�'�s��4��<�|"��eݸ <�6��]��s�s�M{�ʤ��q]�`5qH�j���]��rG�#ç8~��㸛���d+�������W�rj��ć�?���Qh&LG�L���)/�zek22|�l��~BM�q` �9(���j�%Y�7�#m�8&CEVu���TU#�Է���k�P*T8�gX���A�C����`���
n�R���nG��6Mq��4�JX�q��dW��@O���C�7��O�D#��4zԟ7r�]}��H
��r�	a��1RmeE�q^�w��a����|قe����v0>��J��'��(�.0`�{@γ ��L��
�f2�xҽ �qd�?� �-^��?H���x��&�:�/Ȟ<�]J+�̓[�3�D���[3�c~:A��6V�GLm_��v�r�]x~|{=��||ό�C*;�O*���_���DIU�0��6gP�����ar%��π�����9������q*|#�y��<��1����]0j-�f6��$����kA��^��a��y�&2A�Wpޚ�CƼ|�&���mLO> x_U���K <5"�I]Ӥ��{������Z�e��?�q��8���_[� �'}%��.}�����KpCb^��4�xP!�i6��w3ī{'�UVJ3ŵA<n��uo�]s�)v��Û�'2$�rɻ~;Ouh��<��IP�?LZ��'�}s;�1������Cn��s��S�����[�����5������M4������L�9B��l�/4�_W��'-RS��H� ��]4v���c��nL{�_�/��P����=�Ƃ�?[Ї{N ��C�>�����rr�I���+䬵��8ƪ��.,�m"L]Ig�}Ϲ�n��R�(X"�i Q1�������F�ޜ�<qI˒j�9��oH�R)�𱚓\�`�gy�<u�cq����˞��v�o�N1P��,�@��Z�݁���)2k~Y����'0�����8�3y�ZLt�fiKN�)�w�^U����U<���ZK'ȷ`R�RhzY�ۥ:�0��n��(��p����w:)�X�@l�
U2��&��<L`��:@��������>�$́:;b���p��@5*�$�����i*:���QL��M!�l�7@���=C�y�/bQnWۡ�
=�'"�Ί�nnPƋZA뇌^�b���g� ��9~�g��7Na�y*�����2I�v"��_O��V$^�� O�ڞj�Rr_�Y��/�Ľ�{��BBʖ��!ArS����p������ɨ��\յw����D�fnr�'�5)bjK`g�tV�L|n�X���B~)�,!N-��׽�2��G��#D�؛���t ic�$f��V�[M����r��D��4ϸpi��蕳��ě��8D�%u�E|���A��+|�Fد{�Nŧ��`[(IPt��u��7{O�����*G)��"���'8|<���?��ހ����}�+��X#��n�ep��x�e܆E+�t9I7�H��h��R0�����g����t6]^#�P��d����,�����q?8Ť��,�� �^hʖ$�ɖ|`%yUDl�f�.j"�m��`��������X*S�G�a�y#/��azp�4��b�qyؤ*b8���w���b�Ou�Q%K��Z�ɮ軖c_R���J�����$���`c��5���OO� q��D"hg�D6�e[�5]C���ٹԵ�������l��GŏL�������U��U�ɰ�'9OF,�+��!mf�n�\J.��do��>�5&��o�H������o�{���wI����{�*�zؙ]��0��H�w�y�`Q{�I^*/:��\�'��1��G�64���2>�g�����E�2�F.(@��EJ* �B�/�e�t��J�Sb�����ɺ��T��A��J.B�2��,�\1]ᆕUoM��Ѿ�芞&�J��K{~^n�+K�y3�f1kg����akVX0J`	�/�,�[�Zfhu�I���S7�j������g�Q����v5@��F����'���(���V�:�U�nDb8r�\v$A�'�c��\R��M�Z����F|��+�WXں���Sa\Y��4�z��~�0$'����>��ˊNm$D�?���q��䊞��gH��a�S
Es�I7��)I)>7LO�x�KuY�2:O���^�(�����f{����=�b�����;�F��,Á�͇�'�\����W�:�l�T�V�|*7����./�1��1.Δ�"�]���jXl˜��a�m~|������J�_%��n��3��#��N�P�pndӼ�:�yE�*Jx���Arvqx����(������ #!�������s"��-�+sŹ9i�UoR�p��G�&W�+���Մ���O[>Fl?����F���D0#��ѵj ��W��%К�wGo:$@�\�jH����`d0->�'!zP{�6�����{�xR�Y���OT�|_��}��P\�� �b�Ń] 
��&M�'���5DH�/��5����d�����nEE;�FP������֠�j��?���a Tcx=�t(���Q���Y��xu'����ΆA�u�{�89~�^�9n@0>(�/��7�L�19�Wb��.���K��!B�ET�����\ld�Uƅ��Y�`��]�1	S����Q���8�G�Y��n���#3�uZ4�@�0�G2�2M ,_F:��tQţ��B�w��g|�������+}�7e�sE�VN�'�E+�.��Q�U�&�cg�q����yݗ���*�n�����f8�_4K��~��Q�um��q���OJ�P�J��+�);��Y\�����=!�-�m�Tg�R�R���v���ȑ-�Z;���U��GZ��8v<��;���~߅Q������O�(0�tI����v?N�cI3�~/SK'+A��mL��J/G�ޱ��z�� NBD�6���
���������Q^��]���U���߯9J�!0w�T,�9�\
_�)�+'���5,�|4;� 	�vq��P���E���F��|����|�[Qs\�k|�t��SuZ�E��X�����ן�Px���/���
��R�V{*>?�YrBcX%����6.�U1]����ְ���<�'������ͩ��:vS��Rd׸q?q��;�D<˾�{�h���yJ��V�@(jFti>h}g;�̘`\�ή���,��4�&2X�ES��`�*�_�c���6v��k��V����׆1[���ƫ�m�c :�xY�ſa�M<(��At�c��v�6��a��'�����]�(�n/��Eڰ��K%���Q�qv����h+��N��ˈF�i��J<IZH��$u��!����q4����w|XAb����Xtd(5��N�E�x�����o4����C��r�E"1�Vlv���*&ib;�J(�Rb����5X��%	#���[�g?V��c\Aa9Z�##p^%��59��W�;8��Qe�K�ƴS���f����lxM)�y+��OZ�ܒeʼ�'��T7�f���_g1�� /����66>�"Ml��f���̧�,���yPyϐ���%�B����6U��dZY��c�l��䓑Br+�(��T�ⷶ�j�	�Z�jbA�Ոv���)*��a:���@���%!����%�+��]�3�!L�*�
9��6�g���W�y��uQ�J�P�$�	O�2��Ѯ���V������[hL��0O�f�v��s2���#Gv'��S���{��/��T��n�c�8�iz��]�D]Ɠ��s5y�)�\�Ћ=��hm֤�]�`�R4m`ꋤ\�����Ek�@Z�?S]=�X�๲���	B���|�@��,pP��w�Q]�o����n��i&�jr�u8���_�D��
	.�V\,Ȩ�Sؓ>N0+,���ts�씨��Ѵ��.Ȳ&/���g�u!<�����eSLO1l������n��FA���I@|��_ �L�:�����h�,|9U�:6~���jyG��lZ�A|\],�\u^0{��)T%J	���8�7�+R����ז������}�UV3���f�NZ�I�K�d#��X�uL��ߏ����^M���z�B� �@��b��Σ�/�F�1f�,��Ë2%��!_
rz���_��-[ϊ�����C�%.O�}������V����L~VN8c�d�c��rh�����jq�f_���f?�Q9�0�_�a��U__9�5���e�Ŵ�q乷L�F��i��#t�ʫ��}_�~*�{���OQX�Z�[���ڱ�	���=Ⱦ$�=KGL�cR���B0d��
�k� =�Edk�p�[�$�,׬�,�����yh�=�#�[���R�*��\ʼ#�)lp���Ѿ�W�pjA��peY�>Y^�i��TY���0)E�M������Ry�(�p��.	�\��ڢ���t��JO��W�^*���s����-0�&���Qz���������=���V��T�Z�~pI���w�j	qDa�Y��N�0�j�js���A�v���h�P&92�(�v6���)���8��'K��c�������쇂�%�XϙE�͘����2^d,	I�:�,�T�6j�#�+p����v�����1g��N$NpИ�/�>��5P��;q�����'@��8��}�iw��w�~�U���K���e�?2A�v4��1tk "����	T�I�����8z�'�X�l�����@p�yV+&p��%*�?���Wi|!�G��'�e����ݮ��(��\{���Ag�U�p(�8_�@�Ѐ�J��h�}
_ֈ�"JҼ��BG;��z�;<K0逮��?�P��Hj����EѾ��]�-E�\W͹��\9 '&��)�}&V�U�
����f�����wgiӜ����Zm�(��-�
*G�-[��QIE+����쥭��D�_.�45/��;�v�Ҥ�L[�:�
�z�E{��H^��il��0�N0k'�ӶO5���1І�^�K���h�<��m�9D�4G��)x8��7��~�+�9�O˲�$�������W��.�5>eܹ�G�������YJ����xxd\�⺙��E���D�œߩ�����}��m��R�A��Q�}��`-*w�B�u6{�)��w[ {	gx�TD��G���x�b`N¯&����� �GG��V�N�06�"�>-�$�����p
D���߸D�
ߞ�8~x9����OJaΏuB�c&mU�E�����j�� o�h�UOXs] ���Uk���چx*�M|��$	f�MGr�v�5�q�M�r�AI�rl��eJ��s���6b|T�ʄ����]�w�@Sۊ��Q^vT�����T�*��t�5�kO����4h�@9��8N���s�wIjk����^\�ד�b*@R��
\���s�J��Ǌ���4�wPP�я��L��&lGǞJJu�U�67��6�~�N3Mv��_�䵫���c�J!�Y�v.��9CV�쁙9h�Q���$@i���tVD���@grڄn%/�䦙���H�ʐ��~9���eo���:=�8��BR� 	|X�����D�b>#�ʖi1�`��ȁD�,9�f�%�!��I�.اpL�v��|s��ib�'-���I�7z4���O�O������D��9f����y^�QJl�>ξ#/�6ɮko;��s�t����}���.}��6�
�z��"|��K.��=c�f �q8�y�^���(7>��8�A�x C�>�̳B�œ_>ӟ�=��4��r �@�u����4��	cTԼ� ���}���p?g���0���#f��HҼr?wV2�������S]�)�� �2�L�̉b"�Luy��>X0�}�`D�f������xI�"IX<�r�i�k&�ic$: �W�GZ��6�=R��b�Ť9���ϸ��v�6�0��^d|q���s@dyq���T"UJ��#�48�/qy��WW��(��Ǵ��d)�'�j�5qF�F���B�5/ �R��Gu��b-���kʜ�C�ݥ��ߥP�{E��U�!޴5圤�V3�!pD�#�u��R�s�\�֞��)W� ÿ���#�!����0Ȏ/�}�K�<�dT1y!ekf��X���7{�װUg�nN<�id��̍)�;�e����@*%/���#�Yl�����n�+���U��a�*����!�)�#�� 
nǶ���,��(�$KK���'+�x�
�����J%G�n�KHkS&c�!�JW�Z���<
�����4�.ְ�Yg��a�W��':��@G�}�UŦ�j ���[#-�f<�:
��e'W[�R%����ͦ��Z�ʳ� �8=�/g��ƹ��N�m�'ȭ�_)����l����ۥ�Ŷ��ŭ��>��t�L	�v�8<�W&��`�d¨�?��sPMx&K����a;P�I].Hgu���2xY�d�(+��4x^��S�!������R6���+2��
�pB��g>�Y�S�v��WØ�#b*�.k�)=�7kp��)NH��ۡK#j�z@�H���u�;Uր����H�A�E؏o1،r���m���1&m�{���v�N�7;��6=���Y���LSy���%���s4��R��	��jF�#;9,�to�ƺ�Ia��t��}��
��J6���4��Ï�;�rZ���e/D1�����C���I�:�0�J����3��rHUJ�d�z6��0qe?f
W�'2��69�$_]2��":���E��'�=W-��Ѱ������(q(��N	����R
�U�F�ɡ#�7� h؇�jƕn&����FT��*-��"��2"�u�P��F�8ۊ{�%ɽ���\�p�F��2q��(6Y��;��e㈸I-�d?�Ƿ��.���?/�����q�3���[�K?���7�:��-u�ݗ�V�i	�k�`Y����9��Qڊ�%�U�EY�@�mL �؊�����z��-�u�?��:�<��P6/�R�|l���7!h[�Lk�Sa������/"*+��a���!�PO����b$���b�Fe½�1�
8�<[Q�b)[p���{�Jfڜ�����A	��d�a�k�����x�<?x�N�;�oT��ʨ���?WO92�r��4v['a0<�&]w��	��E�qX�b�,=��L����{ ��b���0b*ʬ��}2�ٖ+W�L��Od�g��3�w��:��\�-4�m+\2�����c&<�=�X2���0� �l����6�rR�z��ց�;9;F�mY�s<�\ܲ���������n"�&)� /v�\���A"l���F;&ᣂ�9�r?����d���~��ӅK��d��\~��|z}����;x���\Kl�LB=�"�O����h�u��$SK�����Ⱦh@-F2�3(�7���׋vI�#�ϯ����0&�ea�i����K���ƈl�$^%�0��<��yѲ�+ֵ�����&��U�{U��['�RK�>S��� ���1j���i[��Z�^ +\"��M��~��m�b��%$_�~���Ф�
˭֪��f�9�9�S4�{����5�F�SN&��Ɔ΁ac�Q.�L���.Tӥ�T�(�XW��"�/@k<��[Ͳ���0���A!�tM4�Ty�v�|K��������Z{��^|'+�V(�x�l[@�:�Xrk��9��(�\�m">�04�{��m7�>$�W��[�ٴb���,��'��� �(�T���i� w� m_W�d	"�����@�j���7��9Wl �� �5{�3�95�V��';�a��
����� ��{��>��X� ����RBwC�Y�,�[�1��%��}85mͽT��2�j�bKe	���:y�5���w�EJ��='�g��bn���R�j�K|jf�3�H�jm7�>&�Q��m�R�>N���	�^���z������QT�ˢ2� 	�I�٠T����� ��y�y������o��y��ҏ���s��e��8lM�R�}3�I%R���:kG��`�p�ϣZ���x�[�A̹�/��R(; �]�{ẕ�Œ�1ڢ���UΩ����ԬL��������u.��\�5�Y��h;�,k�0v~�6��|RW�2��q���4$K|f��|��T�h�ɖj;�ɴ1X������)Kɸq���?}��psBM���\���=�E���{鰚Qwz�!���^0�V� �n��y�R��y֐�����I~�[7��@X��L��_�V�Zh��fc�JWc�����k��v4	�[�Sy!4���� M����R"�e���߶iV�ԧS]f6O6"E[���c�xE]�u�v<,8f�;Q#V�r��$�$���Tj�4�wX�i�e�DنZ�V%+s%��}?��P���춐�}oT�`��8�w?M^�,����>&˔�|g���N-��Ls���"�����%W��6~*���z{R��v
��%K+t����%�>�U[HMh�yޘ�H��:�����μ��g���v�Z����G�ۆ�2B��*�̾q3�@����"hʦ;��M8��}�B�������WU�"gf���Y)DځDa�G\�V, -F�]inO8f^���4��'�Z*�0�Ą���Py��Dn:��N��|��hfL5�h�п��Bb�{�(2@m$���,`+q���H���V}"���t�+��̓�l��ۻ�Ҝ����ɶR-^
��X�	7���m�5��l$n��b��t�t ����6�!�k��mmTUD�������6���(��m%ge!�D^���)B�\'3�n*4�~C[#Y����sgͪ:2����k�Ӈ��gBY�cmmhke�!�3]�1�������	5jw�("F��|��tb�T��4��;�"�՟i�=����Zݢ�e}g⛓I�ĩ�6Ď/�8@����?n%!�?~J}$�,�ׂ��gJEn���g8;��-��wθ�'���x �͹Y��)�a��˷��<��J��O_@@19����O2U-]/ז�l�õ�����/�Ff6[3����N��r'Dy6&�9
hn:�`]�z���Mvߑ����*"��"\�K�p!IDk�+W�EV5�/�c1tq�핍wL�);?��;���u����شC�H7�T����]pz�O��"m�����F�?U`ƸҭU�z�.0N4aʬ��B�������W==k9��v.�$bq�뾒&��Z0L��M��fN̸��� �+w�q݇s,���@�l�]�0(Kt֮$�/W�454���sOs[TG��_λC
e��'/\��NO��|��&~�[B+u�
�[�_D�q���/�r��yŴ�Gm�J=͠�(ӈ�1A�p��)Q��`�V&{�%�嬑��l�M~���{�*Æ�w2� |%�Ҏ��=L�Ʀd��l(�9:̃�S'�}c�N�^G:��WQ� �����U�
{����EM�ȑ�Z�8�LZJ�P2�̮+>���:�[�A�y��{XR}��|���M�]A#~'5!A��5^�(�J��h=ַQK���oR�4卨�
qOc�0�2s�tz9k�t~��\��Bi6h�W�)��A�wZ�xu��D�oВ�e��/��_;9�_ڜЖ��	N�����S"0���t�
w-��ЛfO�O1J5I��*�;O\#̾��������I��}!S�z�CnD EK��o��,_�q�LЅc�B�8"-�}u��2�E斍P��·��;���\.�D�9����Сf~2��ڛ7�+ې��3���qz�K�:Ϛk���5L�^�=&=)T�Hҩ ��>�`���ǳ�R�X�
l�Vphg�=��������o�T��+�S	j�1�N�Od2#22o�rf��#��OA�9-*��8��������lWr�fH6<�[?����r#`�� �g	~:��%�i���T��ub��{V[0�a]��S_	�����?*�7"k<(1�4�<����c� �ݛ������-��[���Fd�k
q9�7qC���0[��@fvx�/�F_eZ�sI��j���6��&&�C���'���Ї˟��P�o*{e�E�kF@�9���ٌ=I�7�&E���O�#:�,���(o���e�,$9h���ޠq*�a��cMQ��Sd^���y�N_,%67��I�h@���1�r�@������ix>P׺��u� ��|*|��P�
�S��r���Q$h�jn��]#���T�ߞWS����Z&��v/�!ƅ�Ϻ7m��5�/g�~-�g'P�/�TD��l#͙��N����^�������ވ�p�#�ڕq5�0,>˷�:P/`�\�9rK�X�Ԟ�>�ݫ��o��M+���4c�O"�-v�b!�o����a�Q������~���JH+�-�9�xqM��4������e�H���a�R��W@˫�*_Pi�F����� 'fB�����T��k�������ٌ�m(���p}m��71Y��Q]�	r���i1��]�(�É�է̏���"؝0�p�t�P��4�6E��9�� ��WR���*��ěM�*n�m����#�mi����
	I�o��wd��� !�wV��"��׎�F%16����q��?��5O��$`�˳~7��F~\�Q�����3c���9����
ȁ�cfi�Q7�rTc^�)�������'Hjh"�<�L���q�zQ����k�!�/{��[�~<�7���p���������X���Nxy��5$�¿��ŝ���rֱ���ws�W��r�@�
K"���cV4�W>���6�Yu��>D�|O��z�0_�"�~׶E�ݤ';a{|�����B|�H�j����v)d1yyu�$X�6El�&D�$>ͻ�/��
�#&���?M2������,����%�fB��r���)�<q�����/�:q��B���g9oU���Ƙ��d2���U�)��J#��8F�nj���a������N�"�n��Lda�l#��Q*1��0-�Zg�����1yg��=���%��̞�tYN.�]e.)������t�#��U��y�\�E��=������?{��*�Q�����@��<CRZ-Jk?U{nP�ybR�[��h��X�r+@��*�*�l�ϱzd{
T7��+4�fw�E�cv� �r�\��rn�4�8�|��9�ۈm�I�R{�SRA��W�Ԓ���\�5a�i��>օ<YG�C��������8�� ��y]���0��ߧ�?�e�Qk�����-y����`��ʡ?�����hQ�3��(f����ߨ�%��Y��0��C���}U^("L�Tf�Hz1Labv|�
%��j_1ɔ�W��O�vd��+j�d�ߊWdwX������y�y!�?�%�h�ziW��N���/\[Up�����b��㥅����:�x��#���dS�������� Mx?�p�'�C�.�4>&�b��Ap yi�v/��:��'�����P�e�b�����)�F���3WS�;�Jn{�1&ʹ,9��f\�C{�l�RL��B����_'cb����zjM��)�U��M�?U!^*��I�=�w�95�T&�O\�IN_0Tc��GfҚ�}��M�N�W�Q����[���H�0+��Ϫǚ�1��,���ST֤���-�,:-/�(e�U=[��8�~JV��N�#?���c�-��tC� �� �(�����Y�[�{{�"l���O�-8�e�UE�P�9�ҕ���1X ��8���3��*��K���H�K�v�{���^����PmO_N������>$QN!˨��Xm�q��_���S��O
���d��$m���$j2��y^�.�1�U�����+�|���(�}��ˠEjl������3�Ӱ�0V�YK��#�b�r4w�T'/��S�������x�����+|
k���PO���%ҡa&F)�^_7ِ�m.?�S�?d@EWڵP��I	w1�p���p�*�`���Jx�%�r&$�����b�w�o /��1�c(���1����J�`Ě"�R��:5�8�
�3��Bڌ3��?p��1��k�k�*DT�׃�J&�(ٵ�)s�v8)�����^��v9S�L}�YR.�x�]����VU�ڈ]Zw}:R[�
џc�t�$iہ�䜖����]߸6��KEqj���?Ǣ>��[xď���s5j⡱FF����f��w�7#�C�t�bК!_j}aSr�;�c��������X�Z����u���^�buR������Z�F��R�ס"4���ru�ϥ��H�>�>8ҽ�P��#��2�P��nTS��J�k��J �R�I&�v�ֲ��X����9�*EUb�������'�w��������L����~t����>���\8Q��be򿦢�~�WW���R��_K ��c�����@4���'����r@�<(C�q��9z�Vt���Fw(t�^��8�ֆ��~^"<gw���SPCڣrt���Ym�	�9��Xm����M%j�R��_����s�dX�H�����aJ������/P��>s�k�9_ͷv'S�p�K1���j�vnԍ<A�Z�;٘�Χu-��gQ�?����$j���V��˯�W��6��Cݘ�$/�
����:�_��0L��#&V�m���dɀ�ʅ��|2�գC�/�X������.�Oַ�]��q����3�&j��ڲs�����#�,�ב/����W���>7I��%�t�0�ß�f���A	x��2oP�{���m6��t�sA�ق���&r���\4�`����^�%���̢G%���%(��8�����^�e��l�/��D�>�ڹW�29�(&ƻ\\V��Q����ԝ7�^d�!23n�|�7k_P�h�E ��`Q��a?��W������`�6V�V���8�C���Ҝc>���|��x ��Iv�S�
��Ҁ����3�	���v)Zs�M(��p��7�X1��r����4�:d �c"�y�N�9?K�%=�[*�[L*�ԣ��Y=��E�=E��<����f�q�>���Aoy6�]�~��I+��NǄ�D�{'~�9uD��zc�ku�4OtëZ��}S2��Q�Z�m=�?|�iK������T�;��*�p�$`+��>�o����4�c(x�k:���5���u��b��MX_�`��|��Uw��Ci_'����.A���AfS��j�R�x�^F�[RT��[,_�0I��Yi��[�{<,ǧ?e�S����6f���+Rc����ژ�b�zi�o9+�E��[i�f�����,�BE��dy��x��,X�?��S�7`♄j*,�2������D�|�; nE�ݹUz1'6�8��=���wo
D69�>N4�f�S�ݖ턦H���ƿNO�Rz�LME9T���K��?����=���y ����_��.�)R�Eap��×P���s��a9��ؗȤ��EkYᱞ��7T�@�8�C;��Oj=~O-9i��,�%���G5��cLJ���y[Lm� '�p�0Z����$@���JYN�SX^FH{z9����s��@u�(�۝����y��'���VCL����Uz��A�Q�W��i�e,y�i�o��Y�Յ�"�jɁ��N˺v��t�^�"���DR�����U���h�w �{#��_qU	�M"-�r��� ���F5o�䋓���w�2���'��zqe�JU��k�K�X o���,Hg�H�I
|�ޜ���j1����F��7|�Y�~�'/D9\֣K<E�m�$q'����rS�H�t�\�j�X�~�@n^�k^2?~N:}�8�.���|����<�q�����L׵yy�(��d5RaN-}����&���be��
N�<F�Ј[��V�G���tC���8KM�Y{�]��xZW�o[��O�6ԛ�Ѱǧ#��E494��&Th�ZĖ1a��G�`�;kW��ב�������lO�/�d��.�nҨ(����#^ⱒ�2�9�3|#~�����|t����ǔ�ޮq�� ~A��t@Nl�U�̹�l���Z�$![�g
,VS�[��#�_��Y6�C�x�@%�hHWA�iY7v;�xV9���H79�B� D��T~D����$�s.�Ϥ�k�Kt�V;�V���E��z�=1UN�J�+��� ��:':�>��i��Qϟd�`��8+��ߠq��
Ʈ �7���:i����19^�.X��7P������M�>%3���^dp.��\D�\��|C�]j��.{Y�q�G6���ǳ^*�"�A���|WA	1�pݺ�~Q �OmA:Q�X����Mw�쉶P�V�9��	��ސr����l쭌�(_��-�9 ���z���	\��˔<<\��_��BQ� ��wI� ��5�s�5	}�;M�nն�[���5U>���<sU��4{hԫ&7�|p�������GǙ9j����@�f�����6(k0O��s�X� Z�	��S	�+��9_��h�wtϭ[��o9�E޿A�dl��y u���S<pZ�� ��sn^?s���˃_��ѡ��w-y�'��AK
i�P$ΒF��#��4#W6,$p��_�`u=�|��+�\Q�@9�m?g��[�]��w$�/��Ȉ�\�����ӆ��e����I[��e)`�悻�Xs�t
�7do1���2d^���j�T�A�j��j�sfV�s,��;O�4�\�k'��?=#Ҷ�m!IZ�_��~��H+�Q<�<E* ����ףfN�e��y�[��&��֕u�q\C���b��Iq�}���H���Z��5��;.sU@���DQ����7F��?��B�0��!Uw��	j{S1��6���&��m�y|&�F���9�\��~iV���`�? EB�Q��	Ss<7�i��%̊��9j�)5D�I�M��bk��X���3T��N�L�M{�(NB
��a*�T�$�5�S��M�aAe&�how�{b��>�o�|D�	�����DQSh�zF[��.�1v^}��ɳ���'#9�be[\c��-׫������Dph�}I�.���T&
�*PA�L�6�0��/1��(-�C�5�&�c7(�5{1� 棰�ظa<�\��p�+]}���Ҋ�C������*d�%*�m	 �$��c�n��-��P�T8��u��KICi1�T��IL^z�v�N1K?�:r��#���w,���~[&��D]؈����w��m�/���R]�����Z+ո��D���ݓ�/���d��y��5?B��
?��z�����4�e�[����j�n��]J��놿PX�FԒ2>G���Gr�.��9�����t�F,�G ��oH����i�~�S�R'�1�|�k��p	V�a,�%��B�=�g%�ٓ�/��۬StiO֐� �V�A�e��$���B&��_�RZ�'�y���Z�T��i�q!�7d�8프=6/P �^
N��ø�DqÆT«�cH�9m�̒��`���������!F��"'��]U<�l��l7ې�o�Y!�-+��8�YN�p�h2�R�=EI*������h�]f�73����F �ǁ��o���>���7�.M�	8�f�o�����Ε=��j�a����l��;`���vJ2+@H���@/�1��+
+��i�C.��)Z�{M-p��ANҞ�ŕ�,!���Y���b0�<U�k0"Hu�n�	�]Ͼ-]Ey�uo	+����l!F���<��I�-n������~6i���Bozk�*���G~<$34��Y��',�5$7I\���	'9k���%J�ϺW=y�����O�{�Dr(��'ԣ<��_����ئ����������Ѵ5�l�����3�J� V^�ܿ�\JwF���,�|�x��zy9.��o�w��{�|_��KC�%t��PUG����'�Loeǩ�G�N#�._��.a�2�1ǳ��NC>f���u&�<S7�]�������������D>�@^i4~C)B ���A��j����k֨��H�ŏ6/�$��D��O����S�:H����Qy �L��7j��f�#A��-̩�I�¶��x2�L�)�N�F�4n���/���Dc2���c|�%%:���ND��A�m?�=��Hv*l�������$:A[0uE<���HSb� �x�x�o��-�����	i�9WG3��E�P�:>�ԥ��<�1N�^e�6��U�C��,�3�e}�Z,�Mٸ��V�4>u�:�P4(剡�S�z����+z;�US��V3�`1���<u�b�C&z�i6�\/���F1-}[�M���֧��y	�2N?W����}h�j�x&�ۍM�W���[ZTe�]FgQ�
�Qi�zRͶ����&����n*�!�0�3��yG0�T�G�~I��+�-��K҈X�q��w�l)w�Y��J9S��,��e(<� �;���;��`��gs�n��Y�9m��L�Τ�����}�6�SaQ���c��*��w������g8�j�[����]Q�����[Z��QR�㶄�_�C��k�exƘ�i���
H�e�D���$F�P�9Z��h5>��	��X��֛�Q'������-�wJZ`>�*(l�y _�}w��A��"T(�`
�d,R9���,n�=��f��J����,�w��䟳`�9vBi�>#a�&��!A�,J��􎢂L=y>��SӆK���d�bB�¶�1+��smoK9�W�3a �@�h�š��չ^��y��.m�`�ӯ7�J�'�u6K;{��iN�[�9��E�F��z	��Ua����D���'M�0I/��ݷ�Ôum���.�̞�p�#����#�ޣ*݋vU*���-��z��p�t�T|�?�L��!֐_;RY}z4��H�IMPM��4�?E:��Ԉ��\�j�2V�^t���k��S��œ��ߨ������eO�K�B���>�o&C&y�m|�	zô%#K�Wi�~�o�%z�4N��W�O6=�:)\)���(��]��:��S>�Zd�L_Q,�e���@�Mq�<���ϭ5�E�t�M5;�S�P���o�G?G[ �����H5
֤�S��3�����b�[V�xḄ��N'��7�>�j8���*��7�U	��I@.�^̺T�lko�\ѕ]M����)����`|F��ZW�^�c��c�u�B3\��P:�0a֥�\���[Z�[����?	g䉡lhq�f�|�����2X2��꿟1����^m�ኊ�nN`k��v4��o|]`SV��.�w%�5� ���E?�����
�CҞx�����˽��)��]I7�Ч��\�MVsl�\f���y��%��CD���YȎ�Ž_l�"�Y���$Z�3~��ꢰ&+�~ܬ:���EL�_��ɰ/�E��xVD{ÃŲ+��;��#�H��|���s8���b�&"�	3}=��ff�6k���f �hT{�'�6��:+�����*WĎ�ӣ[��_o� r.����~����>39�����4#Vz7�QI�O�f@���{=PB��<��Z�u��q��^"}�lN�a� �(<z���]�h�&�n�Tw-6�!2	�[e�G�LՃ~�0 �ʊ�6���O�ɥZ�Kn+*e���X+�zu�ә=��	�='6x�dc�}қ\Oa��-JH@KVdr�l$������˟�EoJ��⠒GVM�j��	M_I$|W�OG���k(INӄ,l��C�`��5)
|	�l�r9��h�gܾ:���Z2Q�|z�h!���K+�`he �j�|1�>є}��m��@�>�s��:{DKa��IKO�l�kg]����Af�ف�Z�;�	40SUy��?N�W7q�0&Nē���"�#�b�p%�R�f�I�)�7���9V����sT��C�)��љ��Co�\�Ӿ@�}����B���!�$c�1��D���BY�\�"��Ġ�ʼ�y��$���N�1
=,��X��*�����-^v�u`X� ��5�:�-��Z8න "�*j
{���9��g�&&6�q6l�&X��I��5�>���)����Ș.eukc.�E���=�W=���,֙�W��(����L��jI�!� T"�l^��Y��6�R,*��9�՝��ڳ��
��p�Xh�bT�ʍ3�������R�)=�1/���ޭ�lL-Z竟[�.Ō݃���K���O=!� 1:�9,���^��]��\<L䈫�r������Ӛ�>dv &� |��v��dyX��r�3[@朌��l!�7,a����ړ�廸g�3>pϸ@[���O:�*�j��¸_�ȼ��!ܘ�Vp�IQ���7��L72WA�򀫫2���''};.���{'H&U�*bӲ��N5���O4���|t�a�O+"]�Rg}wH��MO���,dM���w�u���y�b��A���	h��i��[t(*�t����~�����Ne0���>�sd�v�?�+�a��R��%���3��̅UA+�g��>�/�b�"�H��O7�����.Lpɗ=�c|�����
iG,񏦽8����?������.I�C�%�#�*�J\�-W��5ګ���5�T�єv<��lLSA씆���w4�]���g'JT���g�La �c�c��4�يn��ϥ�A�
W����5,kU~1j(	lV��<��N��f��.���~�|P������ޠ�#���zR�:i�G�r�tW_��~����'���/�k)��E�80��Օ��b�)�ǿe�3lk�fcB'3TZ'd
���O���F=Eq:����߈dC��U� ���!��K�WA�I}R���P�B�h�0�����㩞K��%y?��LCFp׊�ԋ6���ל8�]��2��̻���і�����^���Z���՘��o��{�[�FϠVL�eG�q�NZ�,�1�ՓtXW�
:6VQ��]:�go�\Y���D:g��E�������tА!�^{5W�F�?��i0X�������qY8�e��JJ]��)�����4|7	�K���RU����c>/���R�=:�sc�W��|\VFB�S��R���Z09T��%?e�#7{�2A���4�`߬O=��M�\N껢$Q�RȍQ��:��0�q��$O�6�>?�]	<�����_�V#.>L<����V��My?�����;���ʴE��[Ψ��7���
�~ٻ�sW/�yho��@�
���v���%�'ih�>)�4��m�D���g��%��]�,3�k�o�����sS�@����(��VnO��& �4�?D�-��ӧ��|!ܛ�Ύ10�K �k�����z�Uu�h>�=��mW���O����.B�?�59�%�3��O���v"!tx'�*r:Sj�?�ޣ�>n>~k���p^�G�$�S
^ة�z�El��ns���vMf:]��"
�YS�I;9�˔���O�Q\�
z��GX-v�.(����!`c����3U]�5e=h�{�+����Lǒa
��CV܇p�h�ƃ����iH�	�7���<�v�^n�a�9���~zD?�Q�4N��� ��������{�Z���߯υ{�E�����GB�*r�%��� �\^�����������뒵z�<�j�S���H��#r2���5 ki�-���n�m���υ��z�egx��ḻ�3��~0� ��]��h�Qθ��b�/�� ��y�';��t=w�0��qXW��Ҟ��~���n����� #@�G����"V\7��ɖLCmA�YD�d�ߢ��Kr�۴��UJ��d~=lx[H�}���!�<sH���_:5:(0��]Jn����?"r,���ϰ.�v�����3�fC�G�<�A��@��7�1���7���(�>U*�S��.e������?����-�2��+�1洏q^/W��@'Ք�c��0i{pզ��=�л��t����:�A`�y�8�fMg�dq��6}�}���V�+�����X\X��'���� �@�?�ڽ/%����R�]�x�������I�~IR�9f
u�vY_+\)��4 �-<�f)4 x8�ӎgl9S&�|���U=�0��4���%�1e�GLL��6�W���O�
t0I��]D��G��� OLo��޶%W48ܩ'�t}��4�[L�J���!���vՀ%?guo�;e_eC/i/;]���~���{��ο�M8�(�2�l����m��8��4����NJ�(��C��7�2Z��P��C��k�0)��d~]i{ȃ�<U4EZ�s^�A�LVy��%�8����`|�����>�}.��M����*Ԣ���S�[N�/������4V�)�J}���u�z/9B_����l��M(-����g�ҡ�w�͗�[$�h#t|���D	������(ʑp,l�wj���-��Q;���+����/W�2o[�u����^Se.�k�"�ڕ�`2J8�\n��/��=�孮�&�a���FY�&�c=�k�zҥ������!p��,�n�]�Б�4c��	r���;�ڴ��F����rp�������J'�"Z����]�:#G?��
?��h�@�����NEM�h6e�/�Φ |T�6lkXLEyх'kg/[,"�1ZEK���f�Ԛ����}���u6�]I�F�jj���a���+d}�	��bw0�0׊r�/���MN�XM�9�a">�s��ϙ*E�����4��o�����J�t�R��i���^��V���(�Լv�,�&T�tC8\��ц�);�G0�;�\�� �y�
l��Y��1�RX�T�q���q�H�pd�f�����T f�kt`���
9GNx�|3�b�LA)�!���a�	�c��}«	�C?�G].M��e���V~ã����=I���������vr�99�zi���A�FU��#8	'�/�%�d�q�_�����I8���܎�����D�h��5����%w]�k[#�R9�2�Ȯ���$C�ᖿ"��7�y�H
E�� �+e��M�Ήle(�c{n+�5S�!����L�/�F��?��q��Ik��+����� '�mi���
hLjc�#��s3%�����ј���8�֧l�R��#�kDD�[�ԳG���������8�y��EťX�<�=�XL;��^r7�<l�8Ee!z�'lfEFs�/8�������rl����Ϻ��w�H��Pn2����^�1fr�Q�3U��i�λ��e[U�!�JUM��µ�Mu�V�yu����-(AX�K? �PU��J��N�򑪜\�J���ؼ�aX��wA�c�Ii�P���@�-ދU�!cɽo�Lm���ٍje�Ci_�jP�~JR�?���."- 9W<S{�ɜV��,�\�z�ADn㢸��3Paـ�CI��r�]�T�b��������aա�a9�L\Oc�y's��.��=I�vP_�1sV�����'G���Tun;��I�+��]��o
9�/bLѠW
.�T�r3zƲ+��,ր9n�Y�" �(d����4�y?dc�6$�=���f�4��/�*s�J�3Y���{��{B&8���8volxC�o�X��$���y̮_��`%c�.,o�
��OM����]��!�w�Ľ���!l��!\�:R[S����{�L.V\[G_��#X|���: ��Mg��e���v��կn�}����΄4��f ��?�P����̼Q�?�����9�D-��v�"����:��X����A���/���5,4t"|T嶛ߚ��Z�w�$II퓉
��ڸ����~��t�{Ʋ@��W"�xC8�v{h�!�w�����v$����2b��*E��8Ю��T��,֓L�_`�ӓw���иE�B.&a�(��E5����R��c3��7�6S����|� ����J<�٩��~����iBN��T����D�wW-�*�܉�]�\���j��g�Đ�/��T��~WHa�i\�p*�p���L.�� �-�_0Kũ4R�C�^��8�"]���ݰ��jg�%��/�,*Te��QZ��]�
T#(�j�2��2��:��0���u�F�G�XxIq����j]��rgW�}¸���t��f���p���X�N���ᚧt�P�����Ҝ5���{���U�a���B�G`��c�1���Y=��$u�s�N0���̳��U����+���W��
&1��ri�O`�~��B�gf�4���9�L��}z&*X+�+~� ���;�ϰ$[܅Zȝ�ƖXw7��&�0�j\��)�΅t ��/gS�5�Syi��I�7.<�ӑ�u�G�D�i���K�� �~���G�w��ջ�1�0[χ�|��B�5�.�.ya���b�l��o���A��i��R��Kx���e�U���`sI������[������a�s����!͟�5�鶍
1*���ͭX+J�w��s%�#F��+�H�6��	����=6w!�! dL@F!��o�}�+���!�%lJ���?3qg�I ��r��*�HsQ,�Hn�#�k�n;g�݁��ߔ�"��umE�N�Յw1�����ք�m�e�����:e�T:q�r���J�^Y�݆QDU�<�߾S��yL�����L$g|%"�bH�>�������4���۸yq���zU��U`%͠s��u�v)��D���G���l�DC�'�ƣ�������Sk�?�t;��/���A�/Hca���l��K�Ԛ�.่ۚ"�Y	>��������$�)!��K��z�>�X]~`Ep+?e�Y�v����*�=��`����N��s���ߔ�8����#���#,�G��i�>*F�rQ�������k���f�/qq�*�-�6��i&s0��1�Z�R�{O���)5By���1mX����\����v��綜j�?�&o�~�n�	�lU�?�%�����-n�Ohb2�ƱY�xD�9��Շ�R�wy�Y�G���OXί����=;m��H�P-�z#�-�����{���7���K���O��d�$��N#'l�&ziI��2�n���)�f*�v�?1�4τ��������
�|�Տ���	&.Q=a�S�^ۃ&}$�OX#�	��޶�����+Dy�;:��a�ן>�#K��Cgb���M#n�~V��7�;�Dq�?�;���+I��@�>�h�߮�!7�	:�c�ʵ=\+���n�G,ХU�C�օ6%0�>6��z�19Qj�v�ԡQ���� �L��탃���[��}��-�j�j�	R_�^�ԛ~�Eҁ����� 1�i��\��l�I<"L�v��o<�D�,	B��:�=�����f��܋�R��Rh�?y�ؙk�x�6%�Gn���Z:ڂ�����T|
&dr�4�K�w�"ϖ�w@uP�y�C��5��,z��e�{ĝ-�n�� ��:~��D�)2���.�@���Y:�(���J!�%���0��SiΘ���_3���B ���ipp�L�<Ω�OM!�A�4�����K�	���i��3�:m-�ޣ��R�mԕG���B'4�B���0$X�pj�'�b�0��5KE�kh�KT0Aܯs.@�	�1�vi䏗/s�!��ƍ�M'��j�0��j�$}�J2���HA��To�䍾�)۫4�-;8��Y?�(���U����ơQ��ٕ��1��6��L��+m�'���X���R���s����	��(vw�l�6疥�b�a�ԾiѕlJ��-n6���c4h0�V�Jћd��Υt��5���<���Sb1Q{Ԟ�-��AlBo�'m=��Z��+U}����΋[D��2����Ӫ��Ab5ɚJP�����Q�!�z����.	�������9Z����S���PZU��~��C��2+�[���YMh����&����.�s<w�c��Y��3�CIc��������4>)�T�R~lc,�q���Q�V���K%�>���ԋ�?��pr�IeŪ��8U)�8�u�#�J������f[�Ȃ"��"֩�=5W�1�-�6t��!: ��lG��&<��f'�������,�;�Y�F��CR��+s�w9�䈦��	�~�/|���-v�Z�Vfo"��#,q��i3UX;��&�O��'���(ZVv+��㑏R���d�f�*B6ꈾ�ぁ�Q�w�դ2Ke�P��Ѿ�]x�6V���"璜���~�K�[d3����i�16y�h�B�� ��o�6��@���V��I$�i���q�nh��'w�)������!Gm��+��81��>��xv�#��E<Kb�DW��C�>�ANy�je�*7s.eP�;b����K�xH�7��P4'|j7�-#�.) �P�3�$��Vj�&�?L`��g#D��|}
#���I��p`6���eho&$�0�sX�AZک!ܕ*� э�~���0+}�t���"��{YN�=`s����u�{%y�R�Qh��M�Ui9MH��F)�!���aX>�؅+>kL�A$���2^Ю�q��>c���l�.�buahGl�ó,��^�8���%��� ��.�d��ϱk��j5)���F �n�}����#�_k'�~�]S�M�����c�O1�|��8MO�Dh����l���2]��<�\�{k�^�36�J������y���}{62�r�_�Yj��:L! �Ra�[��xIݔ���Ź���y�V��ꓔ�H2{8�����6�X�f������N � ���I^-{��_m���:ƃP��z> ����mF�H?%=��vK�i������C�	�Ը�H�_=��5|�G�����ǒ�"oc�na	e�ֵ�s��CQM��gȣ�}C��$l�ջړ������\{��H��k��m���m�I�t���%���~?~[�L�����sVON��i�>aTn�o���>���5-�2_��r�U��Pl璕�q-������+���y�]�z[M(4}#�L1^Y�Ɉ}��'�j���e݂��E�{�j�'j���G�b�ٽ����[S�q�����q
tb����Ti�P����w�u�^=�&�B�A��`D��|�w���,`s�r&��0ȤSQ&�w�m/v�6P�-���P�l|��)�4�PR�Ӿ\�
�yjYI[�z�A}�k�l=�ز���ػGy��!���k�N��y3|�R��1l�ސfs% K<�����42�ϝ���k�wV��^ڷ?����pwzh�.))Dq��+P���n*Hno�s�2����!�Z��e,)���J�W�*+%*�h�H=J�m�R.N��>�x�E��n˺c2P���)=����/�>�d��Ue�"�����R�h�Q�K6N�6?7έ���D*~�	J��w���DKT��-��a�^�W�*�^��%B:���)~ɖ��f�3� ����F�� ��RB7	ge�1�����Ch@`h)�=8'4���0���z|����(�|�����-�l�S)4�����E{�%��y�
sˠP�& i�v�~B�/����}:��	�po���Zߐ��5��}��s+���Q�� !/��*S�Ҧ��n���f��B����Z>$$=�mbk�-�)(X�rh�lm@ƣt1u2�"����L��E�a��咮�pFs \Ϯ�,[s}b%����2�7��v�RxT>�Ab.Q9��e��ˢQ1�à���$N	�5�20R���䑏2|��`7�Lmx�3�lأR�8:Z�ee�O��GRP:�}����+�� 8���bk��%�>�C��-�bU�y��i��y��P���#&��Gx��@�>�F�X0������j�Z1�[d� /�i� #�0���7�`)�ڌ�vm3�_�U�by{:���X���/��0���1�������p�(�<�́��_/9<��I�NԎ��)L�x�1�!ǒ��"��//!Ѥ:��*m���g!<\���{����BI1:��Ь!��
�`�0	�˝�g��������'E��G���VX��V�i0}S�qd�e��!x��#�E�i��ϰE�������U�F��S�R���@�\D6�kl��8��+�����:�z'Gβ/�e�>o��0�`�'!Qi�:;la�����N�E�%R�Г��� l��P�[��}J`�up��6��F�4�9|(dNfj�����U-���ɍ������N�l�A��h�����<zW�N��n(%�����J���zj�v�ln�=mС�[��T\=�4��FbPZzD�?���q��(�-�8Mp�W5w��Wi�цB���c��H�9p�.ț�����E��	AJ1�k1*DZ:J)S)S�,�TEd���ʁ�s���#=URu�>
)�i�f�q�W�ȵP SO���c|�T�tylu����������z�M� ��N��~3k뢂�Ͷ�(���!H��������Qzb�2ԅ`�W�4����5�Rj<�Ka5қM��c�K�0�f�p�6���P"IБ�/�i�[ŘXO91�?�6m|�ڴ�t!���?�N@V������˗|��7 F=�R~�q|�	/F0(�;�
���v�tSX��!Q����]�7�����E�ZU
mdTx����Z$	ƥC�d� 	=�i�����v;�|(x[���?��qQO�^X{`��{�-sc��	ޖ(���;=D\�X���N��Z뀀�Ϧ;G��r'�8!��!�z��@�]�ڃ��cw�2��E�����iii���ElQ���m=��ִs��j L#��<i~��sQ@Qy*z��Ҙ��G��y���k�C�:C�> o<}�s�|�&��hn��������/\u1E�꒘9�)۟�������������Z]��.��r�Z�����T@X0iy���0�����`�$e�Ԙ��#�68�3�H��%��LiH��_�i}�y�͡Y$�9j�,p�����p[�i����F���������Th�z;b�Ӈ��7�s!�=�i~��@2�p&t��u��_����"�0�q�AIQΆ���ekzx��Ukο0A:�2��m`�\i��B�:ۚ1n��a_�S�I��#�.���yǜ�<8��s嶅�͎q�9tʷ	
�ə)v�;FG��8}l���f�PON7Q���ԜO����������<�]߻��VG��-	vP,�Hi(�.��{�X؋׬��!p��k�lwj��SI��I��|,��W��U�ӧ:���,��.I:�))���ݫ��F�2�dg��娦����S�Sj��#_1Y�3V�P���M@�����Fs�+��g�#��+ے���Sr�j�~�j�<"��j9�od�h�)?�r�>��߽MzЂo5��/�ʂq�Ͽ]��8��JQU�q��
K��3�-H�wFK���*	h��	�^&#ّM0�s������Z�׻ �,Lo���x ��Y�WB�:x�t	�%��ؔ��B%hBO��̰o����uK/~����q�z�`�
�iQϲs���~��~���?�H{ɋrE��E#�D���>~ߡ��i��@�����\�X�1w��xm�+N��G� ��e�ɒ���.���_�%U��|��x�a}�:n?�Sw������a��z"M��楢9��X��fNZ����j�U<�J���¸�.��r6K=h�"��>XrBI�z|Uz������#���Z$B�3A�%cPB�v�W��4�R���4o&.�!��GM�����5���@!9^ċ4�H��OZ)��tܪ���P���QÔ3!�T}�7#��;�t	���G�UF��^2ш?�g��N�*���o�nM�<�U)W#�0P�:�I5��X�O8��#��µ49�v�E�K�+���L�^i�y_�f�}��db�r��)d[U���%@'4�1 ���:�> �N��un�tm�t�j`��
��N�>��y��#$�*X!�ڠ��j��W;�5�0X�g�С�=��n�
^��D큂9��`��J0��!P�(�I�C?G�DN:�!�e�5��Q5���s�i��G_j��^L�
�|��W�f8���{c�hF���ڇ�c=D��RQ�w/&��E9"�g>���&�-$��)��(�t�'��� �E�2���t@Ō얫.�@�Y'lo�/^��xC�zzpdK����d�e�J�]!~�f@��$<�\�TL�~n�d��S�%�(`�W�Ѥ#
"u{�i0Z�!e�q�摌�P��LOK�lp�TvVɾ�N��7��>��K)�@B���*�9������:�Z���Ԏ�����QA$�
�*-)���ξ=�ˌ�aB���\\�G:�`GS�T�.oY�C�~HX��
!�c��{��J��!kQ��L^�qs�g���m+����r��vu�,���m��o�mv�c���'�ێ`Gxg�4F���9����Ę���4�� ݀Aye=Ex�$����Ku�!���)�".��ۓF;<7;�d[wk�2vb���.Cg�e�ELI;���ey���%�'�$��~�|Sݔ0܎�͙�#�?�d��ee�_���ft���
6�L@ZA%p6纵���43Q��;�j�3��R��%6o|����jLPϦ�;��먦�l�ն�u'9#-Y`K������+F�ܖ'����7҆���=;��RSLI�dm����)����e�~�����z��r�ҭ+�>x��/�`oe'�1�ʾJ�>�38w���l_+|�׬�qu��Uʨv0�2%���:=�x V|�P��M�2��yPF`��
�[��( ]E@��˝�H|�'�p~�T��2��TX�[ɥ���^%&'(cd�X�L�诽b���Jr+���x�s��[�kւ#SF0T� ��2���WE���@-�נ q���1�.��;��~aڷ�ϾU:��~���3ggM��������d��/Cj?�����"Na�����x�T��>���6`)W���:����;�X��I<)��Bl�$dף����������n�?Q���j����j�禖D3
E)�|��1$K�>�*��k�`Z2���_��A3P8�;�"pA�hNⓍ{�P�2{���σf�"�ge��|'$�LT��&)��-�{�+��KKیjq5ã��y���ia�d	��J���p��%u�����sX��$��c����j*������Pڵ!�
�� �"�4�ӳ�/Km��r*z�S�~`�=��
U��v�׎�劑ہ�%a�TrԲP,�׉�,j�__/V ku�BwEλlC�JJ��sn^�te��*Y�'�T�X��n��1V|��B����n!�g��X�EH�@�s`��{���&�;�@����kӖ�^(����FO�٠�J�c�|��m��
x�����'��h���q���ɉ�����OC���ϛe�Ձ���;���`Yۼ%\d&��bա�{u��Q9�ʘ���� �)��݆�V;��9�z�))R5iȬ/TKѢԈ��f�ȭ���=c�\�`^�� ��5f����|��3�4!��\X�DH�$Yҁ�k�~��dh�X�F����q���VjZ�smp#2�,5EͰ=�:{���m�87�ӡ?,;��A�E�ۏ ,'裨堘@.GC5��|��0�J{��009*��HeM+�&�#�+S�[���!!R+�΀��X�i�x��o{ݫ�B�6�K����K8����&2�����ށ���b�q܍H��y�_+��c �l��:-��V~�S��>�=lz���{T�,�v�%툖Ӹs��vCy!}�����uC5"������,�Ы%�f�:�ȁ��W��9X�ʦ>:a5r̻����8��󮔍��l�e-]1)c�]���='C9�f�x�F�G���ҝ�)�%��B�����oʉ�� V��z������\��gē���W�)0�b;��q�t9@��f0��<!Q�͐!Qs�9P�-�zO��<�1��,٭�K��p��1P�TCk
������"�7�m?��kW/u@��Mp\��������VU�w�g7��rx�A�G}_��cg�$7U8��[� �Qj��.�Y�KH�岭���K3�hN���}(e��{�+���i�A�Xf
�<���n�2��a�����m>�w7�����FmWD�c���m�0�/ʴ�D�ٌ��'��k?����_^���M����EV9L��8F�ma��o��4t�C��S
Hd�1��/���J���k�ۚ��'�˶�"�5[W�������&�O�5�)|wJ�͠�z�دSı�����ٌC������U[�a��|�7l�K;Dq��EC�F�q q7�}ݲ��2��o7JA���Oo�MRP��A\7��h������!;ah����ܤ�~�)���m`>�r��߳~��v��{˫#�N���Q��������}�"H"@n9.t�i��GW�p��_p�$�o��^����m���s���f��
a�&���gk�	L��"��x����e���~��R���$�е.}yܽC�E�E������Z�9�-�3��9��@��~_4���I0�� �bT�z��a��(�+�q!6Lt�����:��n�69��=ͧh�#��'�͎"ᅀ#�R�Tf���`\���D�_��$W�@�*��r�ќ�zԥ��u�\Z�= %.��e��6�Lғ?������Io�|8P����2p3�u��8�S�߸+D��i�l����?
��E��x��~=��T˭"o�K�"FR�Y;n����Ç�����'�*2�;��mF�DI��w�b�4�����Vu�r�Jc!v���Ǘ@�s"�A�Ñb#���әa��(�?sP�Ь�@�P�+Nb4���$ׄ��٣�u�qKS�9��2�K@�]|`^)5�{����?wO��^��4}��Ԅ���9������sV0�/xݩ*���*����B�F��{Du]P����_�AQ��.�M�b���t��:���6@t���}~x=���d7˥d$W��_��� F�u�fo{q#����\)��2�qZ6���>[I���tZ؃әD��'u4�M�5N��x"S]��"���y �ؔG�YI���S�0�FE�(X;�-�d~N�m�}��X.���|��+K'c/1��qv�5�0� P����d��5\ہ�h�7�Y�j�h�Yvʺnr$�c��8拶�i�jW�ԩ0\
��C�o�I�l�G�TOCR@�ٸ�N�ҥ����$��؂,��
!ثM�Kk2N/�M�>���A}>S��o��k諠��P�zs�ޞT��Z�3?����*�������(�@���G�o��)���T�B��ӣ56����r���Ԑ*�TB��a�v쵛�p��]�k�@�q��DQ�����v�u��i��E(��ÿL�-s_0u$����܆��C3��|�W�}̘�b ^��SZ%��X�Q�k~�cqd�D��O0[�%�@�V"�Y�3��ߎ	]L���#;x)��@�W4�^�R^e2�~]gX���1�z�����[ǅ��%�F�0<�G�̯uCޔA�r����&"�m��t��"�9kq�\�J��LQ�PpZ���a��Ԭ͵an���T��W�p�JgLi���[�D<jK�.=\�?�9�}��� j��,c���M怐�Y�,�Z�0ЏW<��zw���rQ��d��m/@7�%,[��ʵ�&?�8hIS�~���لV�͸��q�����-zuMƍ@]&`}�3*&��t�`嶉�5}1<32���UX4^
X��Tr��A�d��-����~\�)��w2[��V2�v�M=���G�]r@O��@i�����"/�EIu�����"NQ/��e �:Y��RZ��Y�J+�&v钞Y��F��	��oRb�"��x�x�+]�;#[.A�~Q�bK�['3A(4��{3���P�K�=����
�����)���W5���CP=[�[;��I�f��d�k}\��џ����*l/v�18���mC������e�,��;Q���D���~���C�+^\RI��B���'T5�b�0��G��sn����.M�໡�=��]�Ƈq�g�"���~���-��f��3.]��hn��z�B{/,�ڌ ��Ho��Ֆ��NiҴ�N���� >����é[�?�}%U��q���5��d������wC��H�\�W5i&�5���������!,L�	�~�9�<�c�����Ϲ��op*��&2]XE��C�c!�a"xf�!����=}�pS?�Ef\Ѐ�� qG}ci��Hǔ]����ꪕF�Z5����i7J�W��߫iZ־��4w��̈�q4��nQ�%�Y\��������p�CCu߶GZ�x� M�{1_����_���T�XE->�%;$�������Pn[(��8�!`�p
��qRɓ���?�R�΢���]�����B��K�Y����3�o*�O|��9�f	*9�ޖ�*
B�Д���$��<}Y��~��C�W�6q.�"@A����g����i/6ͳ+�p�����(����(��[ Ϗ>$��sE��������K� ,�^2��҃�[�'�p"������F	6��j�o��x�۬�١�Ũ3#�u��X�4?*�L<!��~��qP��0J�Q�m���|��eWb$k��T�n������ϴ�S��������t��k�@�_��~���͹���j��:?B�Ś+�㏮a��e
��U�rU�9U6��)��K{���}y�;��\o�ht�`+�`�t�1�����ʛ4�I�#�������1BT#?I@�<�%9/f-�i��o��ì�k�%������{��${�
7+q��B��wFl�pjG�ϟ��	f~o���9��[�η����uݧ�{�n�I�>�����2VDD��\~q�#S�)La����Lu%�z�`;@�=��o���U�Ğ��(��U�s��a*J�z.���  ��z6Lg7D�b� ���!	Cu�R�����N�O���P�U1v9hg�$��n%�:̧H[�Z�id�pN��.����l�������S���G�����3��&�khcA���d5Xp\)�Qt j�w� [�N�>�����mT���\_�k�)Kɩz7�W*Y0k��2���b]l;���)3t�����"s��fv��b�g����/�ޮ=7t��:	MQ�ϙ�?���)Yv��N(۬�*�/�.؝8].����1����`�cn��	3@�Y����	O����_\!�%넟�[����Ƴ��8sx6ٴ*�E��(�i��g�F��ʖmk��SC}Y��l4+�v���˯Z����\�ّ�ٝI&a��7 �&�!�UǸ]w8����^��.	��ڤ�t����iw��x��IZ�B��4W&�״X��G{���$r�ȑ�`6a{m��i9�;��%Tl�T�o��1MEZ�?��r N�����zڦ�*���L�m���]������t>��	V��2�⋔�����i.��Ϩb��?:��=Dp}صu_�Y^J��PÄ�dW�|E�E`[~>.2_./_�=�CC���y�Cv����d;�CX�㠍�Y�G�cL���r�`Q����F��d|�"�菡6�v��0�Y�#��`h=$�7�"��B����;�h͚0�L9��i�PrW�3�/�E|%gt��?��� hCnmt�v� W�V��� F��	j��Z�d&���p��靶�5�ʣ�=z��дc����׋%��m�M �eq;�d���h>S��%MT�{�D{y�+����Ǯ8C�Þ��昗E�1��|���K�PbK���P5�V�$Q���IkY�B�ӝ�.X���
4�c�As�x|c�_�vS�N(Tf��G�����{b��h{Ԩ�P�1���Qz���qd�w}��
C���X��Y"3�V|`򾛩fC^�0y�G/�핺�p@�?L���,�6��)��M��_ƕ��D8�e��F�i���;7��B�n-5+���pG����;�il��_-�8�X�3��!�ey"8�O�p��e���@���cCc�U���}�_r������B�E�4X�լOa�/�ZP6����@2h풄��78��	����*�9#:~��hZ�[�������?DȬY��T�ޔҰ����i����ڡʐW]"?s7o#%^�,��r�)��!=KK\c�t��؊�ejǗ����_= �� ̮'��P9I�@-�IB�f�^'���U�+�9�'�W������V�_fhutZxVN]�n��e�p�S�:t`/{e�c�N���eSl�mm82>f,h�8�	�<)p���>E�_�L��n��_���J�{`	���;�>�yT�_)B��/l��� �����=���'�T=� �&�\���;��̦*U���5��u�~nw�h]h�P�	�� A�\�7"� K����NwvkU��b0�s���-��囒�����fY	e�|�r������w[L*����VYb�c�7X�K��|�U�*,����!>)w���v��|K��s���o����٦�TΌJՔ��L>��x�ٷǳ�,�-\�/�^OJ�T�+e2+p'j)�W^�֠��?�'�lt9��:�Ul��`�����w�[�����W��M�L?F)\�����?iw!��Zs���\��;ކ^�����ԩ��A�����ɢHx���X*��U/�ǈމ�>���aci�����1�4X둀�M���γ��ZY�=�ˍ�F^^�]���c�N"��Ӂ&����m0���3�K(��CJ���Bg���\�+Q`�։�t�k�7�b%��h�֣���l��>�e������ώ��#���f"I7����/��SYxl�Z�6��rX��|��s%o륞,����.0���'����줋 ��u皟V� �� ����=�z��QZA�bG�t� 	o�hIbR�����\��� �ٗB;�mѲ@W��j�A�B�_Ȕ%�9L�%�-�O��Ec�B�cuPI9ҵ2�+���N�1�KyB��r8�
p��c��.z�P
���8t������Wu�~@��p��S��'ja?!��z�D�i@�HCwu�K~�)x5�1pS⡈*蠆�F�,\�.����[�Jok�(-�Ր4x��t4%�p�������ļ r��9|K���"]4TY�iS�ǭ�܅kXTW�}h)��D/d+Ε�Y�ҿ.ZV(B�j5YD~bĬ
+�G�I�w=4]�7:��YW[״���AR#s��?Ήç�[J�z!#�"� x�vs��3a�����(�AJ���'�V��ef�rVǅ7/�I#)ͪ��e2X�g��d�I཮�Dqwn�ljxq�>"�����;��҂�M!���5����x�F��p܅�".�&��2��c��q�?��g�Y��w���J��cw9�3���A����1��r�4����,j��ڙ�@~���o�?��쟰��V���ҕ24<���6A5�/�&Ct����VAB�~n�U�&9�m.���-��vض>�i��y�u��2x��R��^31�/��R5���4��T݋�j�1�W}*.�D� �Mv��p&�K2>�B���)��%��<gʋ;���c�������$���Ep��g���dq��G�_%��Q9��8����D*T�"�����oUw-z
U�5�q�d���8,��AI����p��4�md�v��:�����]�.���|�o:�!=�o&��O�ox�#|��� B���
��U�-�gGe"5Q�
_(����Ӣ�5^�
&�,�D��	��!�yDP��0�j/�tw��nE��+�1 �!n������@\���77�:D��6�98��~(�EetC�o���GE����et*Y�k.GHN$%��Z4��!�y�������hĲ�*�Ng�Ch��dS�>W~���h�D�}Ȧ��V�~�ꖫa�S��|�җN���9�����0���{EV&F���$�^@���/�@��´1g���]9n�����7��<�yAf'{�g�W�������_�S��R���,������fo�wf&r�Ԙ�'E��L�>���%j�w]���m$�^�w��N���ewU0n.b9�q����t?��
$��V��I璨�gY�Qy�q.Vwr����+�ax�
�="���#�Y��y@����k��_�,�hgꑓ�� �Fa4����_�.c�Άnb�^��x~{2�G���SP][�~h�F�Ǝ�R����rb!���t�W]"��ҫ�{}㭘$��W� �8�X3e���ce�{|�xf/�D+~�b_,:��h��
����$�Q\�0e��ı��q��ޠ+������Ҩޚ��,-P�r�.��u��/;4'T�҂�y*gٲ���d2(2Ȃx����L ����]�I��n���O�%Q�R����y�Q��1��T��w�x@��!+�Ð�o��/D |��-K �G;���E?`B����D+&\$MY�:�t��3b8�ڒ�q�i��O͠������ei��E���Ƌ�hkp�ѧ�ݴ��t;�/�O��wH��4}ْ�F�0�t A��%.'�"鮯r���p�������;:sO�;q���S~}1F��؞�Ȱ�'8�N�����<�{�<���Y݂���خ�U����f�{ƙy����;.>��p�G��w�S��B�h�D��湄��>��q���R��D���O5;�WY�������k>���)�+�?5V�v�ڈ$��)��&e�d��49�@�Gԝ�[�v���[�@��b�۠�=H�Mc�PI;O�2�.>���,�ث�����߮�$|�������K�����P��c��6�Ya���;�I�����h|�(xL����R��	U��_2���P���
�"�_�ʍ�3�FN&��VO��`��U�ԹI��9�V�=��5*�GjA��������y���nV�)��R�ź;���G�R�yB�0D�v��#�x��uU)Oԅ�����р���ufB�]�]n�*tS,Y�(�}3�w��

�/���x<��p=��ƸT��V&�=�AZUs:�xm$ո�"3W!I�_h����+��w ��W�`إz���|)�ۢl�sh�p�������������',Ru����q,4��>MuŠFO�C�����wB��������d �YB_��#�U��G��tH��\���Ӆ�E-o�ӗ�A.�z�������s���"�x��<�X��ex�>�f���M(	oH����}����V�v�ǲ��OZ�ea�H@J�Z�(�1��f���!!��Z���z�h�E^b���D<��Zg9�J.�㹣�p���>���{7�5YaqG�i�R��ӫ����,<��~��-eT���ӂL���bYN\�#�=�~2`��3���t��p��(˙�3��''�%ց3c�k1�3��l'�!�7R�GU̓��i}ʵ]��������E��m�q�e|�N�9k��h�#q�N�~#���R�{�[��xiP�K�i+w�B��r��Y8G<4x�Z�Πf���m�p�pܺ%�w��xL��U7h{ �0#��o��W���޸����T�i�3��^+Nn��Hl< �����\�3�AY��F�6�Kъ7M$�|�$2���wg;�B��kF�52ۻ&����M�'m�v�&��1���nPФ��`΍
j��`g�d�O��TC�4Z6���8X�G���:X�O������ӣ��H4Uwu��S
a=0��P���<g�go%{��U4v4s->@+﷖��lT��O������ޒ應�׉OhX<"}o���we�DQ
�����N��W�8����{�_�T�O����&�/��͊�6xd��[y���1_�Un�rNi�n��ݓ���1�I��������ZDR�<!��;�7�P[��M�U�9k�O�/��q�i�ӇB�ݜd|��dԏ��N�+�#�JgTW��qx�N!�@!]����@(l��"�FCE���?;^B��u���v�y�]�r��z����F-|���1��X9�, ���Fx����;̉T~���թ�Z��W�Z௑�vq;�D���^?@�T`rG/hB�(��U�V��iw�L���d
��v��~Q1�\�]��wV$��D!�\����н�QRܛ�?�?� :_�;
��a	(߅����S��.Ca���W��#����J#����ЏS�fȤ���L
{-��FYc�wy�Y���P�¾*ɩ��>6��8}�]�MOX�x�����N*o4�l�wT�[��6�5$¸�D�Kh�_@��7��)���D���׳��)�P$q-�и�ʱ޵X߼������Fy)߃�j�2�L��M�G^q>0vh�]d�è;�D���\-_G6&�f�e��L������z�z��AYe��1VR)�Esю�����*Ƶ68��&��[V�ܑ&L����ϓɮ�d���3���
�s�~&7_c��qS�����@ ��n�qv�1�d��VK�?��C�a��y��h.�s��W|����-�����b:��)$l?˼�҃Tz��<��Rz����M�#�n���u�b:�W0�����/���cg��X$�H�����+���RXi#�+��y��v�y˦��H�Ne���c���D���I(5��%�dJ�if�|σ/4ƿ������fO� ���W�0T���y�k���^���ߝql(A��X)}�Y�䜜x���B�0!�����A)p��90����\��O"��}��BG̙�˔ve�"���a|����9 �S�5�Г�=�|�e��͘X?�� 	��mv�S�8<EHV+�U
O[�n�`ʨAv7U��Þ���-�_�֯Y��\��HAÿ47��8�4�߽�[�Χ�l�턠R5/��`+�U7T����4�ZQW���.���s)e��:���;�Xʽh�ܞS�?����k٤}֯�M�J���=��6v�蛐I�Ǳgn.�3�N%�p�o�ܙh0c���.����z���i(� ��m�_zgA6<���4N�;�?��O�.���LjrZ��oc�I��XE�Xw�e�D�_��TX��x�:	[ē����'�+d�3W��DJTT�%�^�f��L*[��~�U[����Z����bwo�Qw�<`X�����0����f��q��{6�5�ސ�8�`'J��Y��x�&�\���m�cn�P��^�Чq7u��z�Π�	n��2i0���i��;�"��wn��t�*��5a��(eU��g�Ҫ�mU)h`OfWyPA{�-��ŧ8����y�%	�\M���X�(
�ﲧ)&���.��Bg��8ʴM*�cu���j��̔�M~��P�X¦��O���	��*��T��7�@,�T~�hy܉���	�yE�h�<e
��ܜ��Os��q�5��h�Ve��� >j!j�\d���5&v5��%5��~��aHy���Tf���vm���G.��8_�-�A�Xʐ�مlL$��Y��/����
�h�u�U���=��f���V�@!P�K�y_x�C&�p��g<��B�&��OӔ˥�u�Im��נe�}�Z���'C��\�0�� ���dHN8���Z˛;m�&�L#��¹�	U�����9cO����'Ș�r������\��$�I��Ñ@{ɭ	,�~"����rP<�3~]��X�	�� K��g�,���e����R�W��E�̱9I�tA�Ӄ�uW�/��g�R�6��J��ܯw��%6��n�ϯN�J����m�0�8d ���s-�!��	o�vF����%j�1��L�Ye%w���=J�ًRo��wl[�Fw.�MAT�64�7�4PB�@�yR	���i�����~��5Y8���
]��`��#語���h&��Ȳ�(g�<=��=9?�/�H�F*X��K�.�<$p�ZUy&��K����ڿ7sV��A6.1W^6�=ު�z|p�C��P��AU��i �OC&Q��꺴3C�(l?�g�ɲAs8������1z��sᐵ�(�hg`�0�.ENL�;��eSă���6Z�7~���W�/ϋ���z��i��i�Ś��x_9��v���Dɕo�o����&�;��RU�n���G����B�2��x���<2G]_�[� �yTvR��[*� LO�+xB�ɪk�.�&$ΐ�o���ԕ2* {6�:��L�h�rV��8���k�R(��?�M�x�1���`δ�j}�c��:�Qd92�/]W�Bn*kx�R_�rlɒ�����HU�7pڧy��5#�gP��-c$�?�ECj�-N�e� �(+��H�~��˛?Y����5���#~ƙ���R���4�y;;��yh�r���(�z��.xp�%�<�ޠ���9�"DT��D�:`xG0/-�Dd��ą+�֖�ֻp4�o(Q(4���a@�x}�&�n���)+�CnaL��_vi���|��.y�"�>��	�{����X���& ���S�D1�����OmN�#P�
����j�0[ʵ8�Gt���hV�Ŗ
C���3S4s}����oJoZ|�U���C=����h�d?�#�D|b8�A!G���t���@SJ����l*�Gi�'��l$\��m�T2����n�9h�o�*]W�����E�D|&Ļ�l��c��W��<���i��'�����3+�JE�p6�Dl�d����+R��_G�p����ϵ�I��t��]��x���c���xb)VM��Ú���1j?������s���W�Q���LL�m�;ΠZ��"��Fr��a��^����br,MV��Ӡ`�,޶������	eOW���
0z�����jw-AL��	�ݘ�t�%!j��γ[~���a�bJR��ѓ_
�q7���������⺸��4�i�D�+�47��Bt����������ؠ�,�.�KW�u5����k�
��2� �-c�����Τ��6s�o�v�}Gw�9����c�Y��y��j�H�m易�$��	��A����a�l[�2�f�M����%:�浀��%m�[0+I-:`-}�\L,���d�m����vV</ ��LN1�uΦoU:nE���.!F~�i����u��-��?�K����?/���;RjU*>η�����VB \����ʣ%�ۀP����F��<X��z$��F�|��mE�"���f����>�c���w��y1�7�����f�"�'��@�G��O���� E�(��?��g�'5���<f�^�@��`�:�������_�vV�D4��"��~Z����Qz����h�2�"�L1]�0ݝ��Dx��O��ǦN���U��%�6dd�$�-~�┐�����kr��"<����`������%"ic�8�_���타6#IDX�d�)W�~*�z��_>U"�e̎�!�EĘr��Ba2�/�4%[j�B��g��~
g��Z��2��	7��,9�Z �p�����$�ǅ���у�[+E��S�EnG^�Ϙ���p�Η��>�{1/e�}�f�����B�� ��;��ekϧ�0 ;�P;��#7�0��r1�v�U-7�g����[y�lR/��˵�V���߁�xp���ⶮ���py�{|�W?���B�m�"/YX>o2B`������R��'l�w���t�E���t��0���k�Ê��{�&W$Թ�y�O��A}���A�~j���V��Mם6��I��n22H��e�����ǿb.axΡ�*��_��8� �Bo+��6��}P^D8n>&9}{��qb��o���߃|��K�ڭ�B���w^�z�~���N�����5�O۾F�UG�~[K���I�x�|��^�I���>4^B�n��*i��{�`�9���f���Ua����!oU�U�N��6JYnP���H�+
m8ۈL�bdX�ӈ5���E��ۛ7��*�e�Q�ګ!cu�\�_^�����Պ��y�_�\�x�,]��ٱp�_�`�A��0�;��|Y��K��	��h���NA����(@$�J"����sл q���	Mcr!@��,���������N�	��:ؓt��8���\�8�H#[��!c�@,�z�u1�n�I��VA7�~@K&,� 1 �Ǧ�I�a�t�#���{�:u����U�6�2gAݣ]|X�hg���$�ʩnt�^���mi��3Q�z�y�#�|EO�Ry�vz��O�:�@e��3Ğ�uK��c{҂hϠH�5;�<���3*^_�z�J��v ��x�����k�����˴�#=��ŸɌ��h�4��U�	k��i{�SG�7n�[�aMId$�J�E*����}?H>�ο�P�u�P*J-h~��s��J�V6���N$�puOA��}�[/c-���;}~�ˎ�m$���s�N�u�㔁��͑��9P[׳����jc�����>��s4|0� �����S��~K*�tF%F2�=,�� Wӫ��ީ�������rr��|�daXVZxD���h�X}ز�{i}�F��{���0������͚�]3Hrc��s�0'�w�t`h�����U4*9���+U�B��@�-S������.
�`�p5�L��ߎ�/R1������W_D�#j9?�1�V�*2!����bv�>htg�ޭ�t�E�gas`�n�WP~�*����B��_��z��"��I𫳴W��45i_I���<P�6C�cR��@Ș���ӭ���̘��
Q���Rᖉ��d� ��P8��p�O�h6x��� �������F��G��"�H�i�n
���;���&O\��mvV*��f��G	�.�į��,�ͫ�ծ�ő��>ǽ�D��w����o��4��2�������>�p����$���gQ��j�1RS~ݳ�#�Fc;	�׻?��P�[B�9B���5�Y/ϐ�V�+��2��1��Zo
�Z4��h�tԲL$����;�<[�X�R����*ꃒ̀���$�}tMD�p�Q-�,�h}��f���y�}��㊿�[1�::ӧ#��,�
\!�2�F,�Q��}�]1	7�@��g�9���D!� ���}a��eCc�((OK��tv����a��H�W��A���n�a�4�տ���*<n��[j.�H���T�����f��!�snVu���ޘɗy�8^��u�G�ȋj�
m������`<�'����S�x�*֩�T`_E�/t��k}���Lā�˓`��L¡Z����e�B#�B�p�h�P����@�h`~"� ����Y�-������}V��r���neў�ŉ92(��H���T�s�E��R�V�b3L�G�K�t6��#	: i.��6�����a6��Z�I�ih�<�?B���t�i����'��æ"���ƌ7y� �-��Q��NvV���
1�x:E���1�L����-����X�i�K�z�5��8׸�?�Gc�X���js
q��	�B�'\s��6��ts:�ELI��gԵ.��Jz	2���M�Iɇ��S{�+<�����Q�g��j3J"��R��Z�z��@[m�������p�F�T�u���wՆ>�Ї��J6DP�t�m�S�q��b+e�ה�
�hǶh���P��	?�� �-A�M�e�ה����>��3���c"4V
vf�B��Y�p��]���;��>E�+Z�f�!#$.\�;�H��
fڊ����m�2N�p�[~A���NW��^��Z��%���W�b~�'$��)l^GO%�Qo��4/�"��
?�6ՊՒ�l��H�����2�ժ��(��t��|�=8��{��ygf\�5d��$Km�Op�V��`xXyJXy��_9-,��I��4�������̝�/�m&Ρܜ˱J���0���(�KT�5sh�E���<{P�vL�'vW���j˥U �2;*(ooP�}@^J������)c��r���\ʲ�Q���X��	�0J��
�O$"�}�I��5_��tD�Z[�Iф��5���:������-s_+F���	sT6+)�׽�J:@���;:d��!K�ܡ�����y�8cY��¨���RA����c �� ��	::+���i�G�e�F?�}�϶�w�@K�~�	I՝ېC��iv�L�Ia��S��V@�]��qS�9tf+��\�i�{�*��Pc]�����8]��t�Li���<%�g��
��}�Y�J��7D!{ �u���Iu8�h)'U��0�F�RF�+"`޷����T!���a�[�d�Za�y��0�ĺ8�	
a�vH�������S'�zS���[7��U�#�s��a5v �D�18b�K$t\̫*�>S�/إ)
����
Ug�;���P�����B,�=�"W&�t��3ѷJ`�= v����]�2��G�ݚu����e�8(!+(k7�����`�Ld��BUPX?"��~�T����T��Q۰�]&3G��BU���v��B�\u�+�9��q+cҎ�����o�<�Ѳa����� h��z��G:j(P9ڋ����+�T��� ��]���~6���:]_e�Eδ���1U�=f��P���tźJ�گD-���7lL�ִ��Ha�YE��iZ�TЦH��-�7��/I�y�+ݩaQ�l�Q��s��|f��Q��T"�I�B���ɦ��Rw���ؼ{��rxw"hE�=�ɝ?0@B3�>F�}�!85��r�=!�)�����䱜u����[9(��=��1zl�&N��}���ȿ.�����㟷�+M�����<��u��6�`KbC:�;Qۅ��aG�ʹT����:*���_��Z���6�+7���Z%<��|�[y����%�@���:����a��F�gj�����`a��w��0�@v��Ԩ������g'ܟ����ؚȯ4����@Ѩ�w&��#�9D�α�̪�.K}�@PN��>^s�3���8S�C�K�����ǆ�}�$��� �Vvx5��H� ��po�g���|+���v-sԪ��"!�e���ݭ����"�7o��!�q[D��Ml������E��r^�%!���	��h�uoܱ#����'+cs�Q��h�/���������hh��L�Nݹ�+�~{����b��c������oc�-GPi}�ݧt�	�&P]HS \ߎAw��$�E�]�9��A ����{���)�?�;+�^V`Ӿ�(�("��_����nL���?��p���9�«r��62��u��C�Dڑ���^��F4ӇEg�ܬ.�:��A{q��t�/\T�V�K�ݲ���;�7�l4��S�/;�dX�^���'���Dh'rCO=�qP��'5u����?�"�5���'x���0ݎ��#[m���$Pޑ���(��"h��VO3s�R"J��^H�k�y�+�6�l�&c��|;�6�?y�����D>T������^� 
�8��o�\�ֽ�щ���W�<Oʒ�����mA~����zH&L��zK�����!?gpFTT���$�9Y��Bɐā�5�G���r���K���ns'8��Yٓ��h�׹�#\��B#(v[���ڹ�G�i�W������H�F�XPNy�c�̎ҟ%Ŷ!���R�Unr����l��ɮ��u���X�1eF�2��נX��؃[�A����
�B|q�$ʡ�K5��#�#��:����O��Ғ��i�Ib���"��j��%t��٭K�'�K�Re}$Q%��rS�ta��E��Z�f;K{�mtEVd�	j1�jב��q�j��>��/��z�uk3��59�P��2]¬��������7*8V�z������Ϙc �/?�P�^ԃ�+La����!	�+���g+�BHѪ=�#Km$���l9����������~Zv�²��淪��@��.l�x>h$��y���<��x	�ӽV	��z�,'�ذ��[�([�����N[�\���t�0���t�o��~ߧ�I<!U�(�cBK{�ZB�N,��r�m{��W�c������$����|��?�ꖎ���TVgU¯}��U�����m4�.v�����J�}���	Tԧx�1���I�q���k����C�Н8f%���@3�_h�EU�-=
�n�p���i����T�DQ\݅�|� 4�U�E����+�-4�P����(��X���-��zT�Z���i�d��\��)oWk�+��o,Ø�*�=ܦ]�ۓ�,\	�oΔ�]<^�&�|��(0 yQ�XV]�0����4b��S9o;Q��wmFZ�y��	w���☠Ë���鵕נ��ьG��e_G4�!��[�>��;J�Oq<܂M�gv��»���3�22u6�}4p��>pR]��_Q}�4�w�B2@Ivr)�0Ppa�:�����kf��t�C���ؠ	����[�b�\8��4��H��VV���[k�ϲ���A�x��]�η�K�ߣ���&����� Z<��{��-j&!�_��˟��NE���c����m`C�X,��\�Zj"�����|5�'����6]�fo�'d>�������U�u���K�*�Xt��D��{�I����ɧդ�@�$�Fqk����.�0<P����������Y�?�o�ɗ�n�$����MR{���H�Lg�(�D��.D;� t2 �۪�WZ���ʊ�7����"~��-ۊ�7x b���t�_�e� N�m� �e$hIIG��e�x� �'ICHA�"��`	'Ð�-W��;'`�w1�Hj fv �(	���E����kc��ۏ��f��޼sNt��Y爀`W��@��4�����6�l�����5&n���A�֩(�%�E��|U�O%��9��K��WoN�(�kX((Z�Z/%_	��=}PSpE�����[���U��� 2,$/`K�X��`EE���k -��P9ǻ���q��q��uѯ(���M����B�a�3{�D�-n`�X��XW��5X֥%�2�HI��.�(V�U͛��)�ދ�\�ǻ��ט����m��؊x!��s�Tg�i�}Mb�#�nLP���bAK�'�㖝�FM��x����<K~0m[�/Y�A���5}�o�%z�-(�j8���m���L�p(Ig��<�eN��O�{B�����9���`�1Z)����_'ˍ�B��u���\�?6\��) i��QIv3�����h�_�{�p>V�#�4%U������h��ˢ]'dx�)�OVA�z���dۙ��Ɇ�&q{�I��;M?���ʱt�p�Gf�����?�kZ�,�|L��*�DE�5S��?bʶ3�8\ t�+I�
��6���ę��.
㡌T4�)���F��*�:.�7�n�j��/�}:X�vỏ̹�' G�P�TP��"l��ۋ��s�T60M:%�Ye����K�!MC?n:g]7� ]%�=��d���@���̊�F!�7*b�W4��EObS�	d�܃i܏��J޿�PtJ��h�ջ]D�r�u��,�4G�!x$z�����kMvnHl��D��M#_T�,iI���/q�ǡߎ��
�dIM4g�T�P�k4 3�a ��/�1�kVh�S��r�̡UtT;YR���9�}�d���Tx�XB��[��A�6K2�.��g�7�{�[����;[���]�=Z�$`D`~��}�����[�C�Y�e�S�K�)��2R���{~��Z	�g_�Y�X�$EH��D�K�5�_?z�R�n��Ê��������|�����!&~��kzI���x��PE��^�ǋ�l:%,ӺE��˚e�&8����Iqo��2�N�lf{S*_�3���ֵ����Q6��"��������\_K����T"ֹ ζ���*t�\�m�+^�n=��^%e�z��P�aPǃn��:������T�DD������$�5�ũ��O��L���L"�C�/w�zh1	��i[��s�f�����?ɋ����k_E��2��櫈�a"�b:`�r'h^�wוdx��7�W�D^v��騘�3��Fo�z �&4SzK�Xu��(�x��"���F��} ;k�[B ��V���~D����>@%���t�}V�/�
�gn�[�V��e���B��4>yZ$H[�%�F>�x��Ƕg��L�ߓZ�׮ꖆ�&�0�S�g�0,G{	�,������b���[��;1��������Fl�����p�-P������'ח�t��R<u��2X���{�NG�W���D�]r�V�rH>�tW|���>�"l�f�dgA��4����w.��$Ē�}f]f�!���~~�L9&E^Z�ԕ�P�Mrx��&����iK#��R'��I�;��a���ܢ "h�:2qz؂�&Ob�r;�R�j�[�-�T����OD�Ԁ���֋��k�ޚ��p�)�A;���:$�Xd�|�"�&u?&6�r?���9�u��Y_�|�l@�*�\a٦�_
~3�lEs�X�r��y�n%
�o�������3��dz�5���K��
TOi�ۣ�ʧl�X��\���lx��
�4_���d�/�T'q�M��>�5а�9Å	�H2�����/b��	���Y�A/B�d�T��9ͻ��Ǽ��O�"2l�!�,��qv�|�Kc�@m�ح�I��,[��Y&�P�w�*� �������ʒ��k����&��B^1P�F�o����J���MN%9����l��I��w4��M�7i���"����%H�)��=�r	$?�fdb}��-\�\�N3�;��1���C* �� �g�0����ȇd�n���I����[��{�	����%�]�9K��ݗHv���i�Ԛ!�(�ߦ����G�tZOo���ƛ߃lV�;����ê�;�6��{2���H�
~@�a!K�,��C�F��<��N�5�������xg��P�"�Ar�کJ�,��\#A����w�͎�|)�>��/4!��Ƿ�8=C�$Hd�	����fK	G��k��4�$U�i�
H�3>x�%�J�M׸_�`�c�Dw�=�O�j���vl�Zp��]=0:o�*��k+v�s���G�1^�c�l'��0��%��K��C�X^�!�G����UV�K�O��HMh�ٸ��_��n,������Î?�?XvT�W�-1E�F�k	�Fa ��b����ڱN..��M�/Zwa=A���u�uz���!�<�{{�2ƣ�w��d����VN��w�[.�1՗,��sGԓ�5��`]z�W��J��D�^�8�1�/"b"��fp��a�$(��	�)� ���M'��Π���J�ߥ��22u;­նz)��~��ծ��u�L!�[����lҾIrٶU��$W8f�șI@f��8�?����ʵ�t���Y�x'x�-`!u�V_Ė8u"5��۞�:�_�E�=��P���AFd���+�[���k� T��H����V�]>��/�n�eĂ�,��V�"f;$.��s~�D�k�AS�H@��J�a�9О5�.�w�~��s��йQ�"Sm��ǚT�w�����wz�ʦ¹dE)��A8Ƞ�4�D�r@�Wk�������	u�8��a�B�=ߊ�ե���pef���Eu�m�y����q?.���в`�ZoF�7�J*���c6�b�n.�.7fF��G��-���������Ŕ��Y#�k�&B^U]��������d �b/۲ec!�hkV�J}�|�����|�[���X��ǌ�Q9E��0E��ҧͳ³�����\۱��!�rM�-ġi��[힬@w�����gG�/��[�q�փed\��Ӱ5�%O����Me ]y�o�o�^ �u6�$�>K��v��Cю/��˿1�h6��̩�K�kF�����3�/�-��ޜ�M5|�{!g���HJ�����2���9����wt?��G����s��R�  ����k���!yq�9 �h��8��ۙ��=|�.L�k 0s�z��8�W��tV���a�����*�{����B��MԖ�/"�U��C^����Zkv[���V�u� �����∽�
�U�A�lLX
�/ٰ`��*��װׅ`�4��iG=�oGq���w׼�'�}'�p�_ܟQ���m�%UDwm�q��Z/��?ȩ��9�ۯ5o��� L��cܦX�q<\�O�2O�yB#+��oIa�����l�23L��|����3o An88�|$�|��R�k�:L�bg� kخ%�"E-�ω�b�]0L {�9X��]ghB���Ij݌ǆ/:+U�h�DU	�����l�P�LN��>�T���6��J���(f�{�]R3,1�{�5+,k[�0q"	��%gH2v�Or�Ԣ��AX�\Z�l�EeǦM"��.��"���*g˛�E�
2��.�rn۱@��`��0��I�Wq�j�I7��8V��_�:�;�����b�W�ǥ7�JҜ�i#JH�9C��+V���ʘ��s����M�O$��{��K�
�n�5mKsXD)4����}�2r�� �5�HTt�n��y�u�Y�,�šH&��;P��.�,̗�Aa$��#�.��E��6�y�dC��F�;�Km�PF�f��z�6o^�P�A��A�3
7.O��j�'�͙��+HF�n�0����`:ȍ.`�bl�B�9�NQK�/�it^%�&硉3<ػj"��Qi�����E�	����k���D������htM�E�P�DO^P��̒��r��x�ʰ>|���8,t� 4E��.�4��߁�-A�54sXmP.�eg�y�G�br�OZ�� ��Ѽ>\{ҥ�tq�œ�@wx�v�l�I��p׊�����*�����u��%��7O%9�2���rO��ܜ	V�G�����X#=-{�w�L�Az���uj��}f)�!�y_�(�k�e;�.Є�BG�q8.��%�
��B"��	#y
⋈�<(s8����K�Sg�w���/^z
W��g6Wq7�!�m����E
t�ǖL&�Fi
 '��OB�
���`SΪ[rR���#�A���ΒI����Ζ�_]�A�zu�+1��O��<M��Q�N��Fw�IFھ[.*�L1�L=5��:jc��nb&����G���|F��A������T�KU�CI9�+ &�B��J�%5#z"ō�n7�'�#㉆��S0YG	*3��P����fUyUkG���I4,M�����V��VB�p���sE�*���*#ٮCҡ�,�hAfcZ#��bX������R)�w��T�*�4���;�D,i.�L)���_���eK�w-�_�e�LK��P��V��ȗo�g�<��<�<��]��뽂��S�����,)AzxDГ�
�������;k��g��*�D�������<[�J�lo��[k�By��o�u��3��W�a��aO��y�4�cz�B-����
{��(��7LVD�S�i�޼-���럟b���2� ����6��s�ۊ�i<ܼx��F���(���"9��������E�#�u��'-� �nlRtzm҂�16F9W}��F�Q?�Bbދ�[cɽ�Ut�\���MI�üp�����i��KM����V����L�Q�Sg�q3f6.����y2��@ę,c��Fp��^���]�<���{u��}�Q�Fid���ĸ]j~y�Y�������;�%`��D{�|�e��P�8��:"��"��%)��YX�)���������Г@������˲R�sIq,�^}QXm� �Vo���� �1�۝��*���f�_��x�m^yL�ӎ������:rО#�����g��b{��KA�54�#d�dH=�;����RJ9�k��d�3�$Ht��P`śQ�+����v�����x
^��E܎�ລ��%d�����D̳ܹ��g�׵�^�X�H��XzgózEԜn=�4;����і�/���u�?%���Yrb���92z�Ժ�E���5�"���A����S�J�l$��n��;�Z��/8?Kb��2S�9�0!l-�8����5�OB1N�x^�+�@�}�]Q�^��#��gsd`�����lk���䠴1���)�!;�Y3L#��N7(���b�]oi4.��?k�e4��K���!2x^�4=�	'� ��3J�t]�r��q9�(c�K*K�X!?��Q��ʶ�aq�@ƾZ���pw䩇k��i���#<r�ʍ�o�(�M[�T[���mE��?�̱Lp�E���U�	����A+�Q*0��wX��4s'C�Э§IWu�r����7����TbGC�Ɨ�ꪒdY����zH�u�!Xd�V�Xs�s��~�dܞ����9~��y�L�Y��TsqoI�K�=]�Dd�����܆U���E����ϸEUp���a��R���,P}�Blr�@Tb����>�NT����ϋ��^�~^�F9IZ}�O��t�!���i�$�[�����=�>?�Q9�C}��.�*M�3�gn$��s�7������?
MO��_��ځ��� ����oE"���]�s�I7/Q���ƶ�IB��+`���,P���N����xZqf�vd�3sN�t��11Yy�>�ѵ�c��1�n���&T��A�R{4/\�eA���E'#�k�8p�j�O�=�8�^�<A�l<�(u!�p�,Y�� �VK'���x����&��ږ\Ų
�9�+|�����,&�8��>&���v6E������KQ�/�5I�v O�Gʐ�+n�)97�67���"Τ<x�ßl%���-�����Ɂ0���2�>�3ԗ�&�ݫ��bI��OQ	ZR5��È�������YT�@�����F��b ,[d*C��5����(�M+pS&
_H�\�k�`_T���0U_ܯD����hY���1�#)�;'�=���nӋ8��j�^R����b�h�?��N]9imF����d0��X�InV�FAP��6R f6Rb\o�)e(�3�������u��O�ԁ+�6%dc�PFY���|����
ؾ�� ��ʥ6r
�U�N���/:�J_��0��g�����3j����ߋ8���D��7��01�R�m�ȹ��ye�rz�˩���=���֥��&E�>-�@K>�m���5jCP�1!;Y�w�R���X�@h�����
��d��s�&w�n|�t�S1RTd�u��	{q�I�� �&������ޥQ�k���$yB�O��W{V������DJl��K���(�o:�۫��ɟ�� s�sT�6ƹ[˕%L��Ç+b(z�|�Mh��%��"�<�zY)�"�R_zp~��,#�XbA G�g�21�����ߠ��,c"���g���<��mqp��k%K�%��)�x�a�N�����Q���Z1�Eu̱}N��*6��b���Ɨh��QWy����{�Q�@�BP�O�����R�2�X��*�����ӓ�� �)=~\B�!3t�rfٓ�c�@
��w�4��|p$��N��|=H�f�Q�c�K���9����p�y��x��͐��C���k?�+&�ǟ���Bۺ�w0�e�����m�R��wg*�\��.�SK��� ec���޺��S�o9m�<`<p�ʍ ��A��@�7����!׾~�S���3�:�Z�7�hu�_9 K��8Oa-\��
@T�AѭCƣ�>jL���!U�&���#�%���1X��-��t8�7�jpf��΋G��ʉ鶵U��X��N:�/���/�IX�� QF��� v*��¾A|:Գ�c��ֿY|6�H��/�'�{&�z��<Z���v�b]C���!�:�'F���<�AJ,�FC����lVrA��$���k��p���1�����HC{kl��(ݯ�loA�1�O�Q�����j�
�n=��cc�m+M����ѧބv��]��ʗm���7�ì_���bn؜>�}����*�_�:�� �j_�$����ܶ}�?y'�'�n��\G��x֣-����u\p#����4�w����vȂ0'��d�AV]wn�"����?�N������0a>�ܧ��[W.���`���Y�L�Nã��8�pA1U��B��>���K�bt��s\��*�-7J��1�E~�7�7R!��3鹯Į��$1�5���G�,1J:�Ĩ>ɰ���\��,O��c�J�o�c����k[a<\7�b<[�}S��.W^���6��4z��"o�e�d�E���8<չ��3��Y���	U�j�C� ��Z�4~����I{��Mܜ��g�q��(���l0��UP�f�M9�vOW��;��K}�����#>���B��v,i����� ���{��Y��.Ɨ|���Χ�꼥oG5G�f�
8�Ã�oU�9(k)���j8͓��	�r�K`������EWP,)���2I��Y� ��!ĝ+��{a�� c8;1Q�?!k��� ��Q�)�a�wԓ�ʛ�5�1&M��L�1J<��\ݟ)c�,Ƕ������(����N����a����M�`�~ek� ��F�">���	Kh�<�_L>�q0�ِڐ"������e�-�iZN�*�[L�%]���9	)�y�	'�Xq�a�>ƥ�:�0%�����of���>/+8Q�F�e4���~�B����Y�+�)3�8�|�k�UN׏��u�P��&e�v�np �:�jy�~�З�g�趘jJFo�������?4�	���@���#( �w���1�!������Nބ�k�8h/E�52�#��a�:kO���o\��C�nS�՝"��*2�fo*ʅ�ף�V�R%������Mǁ�%��F6z}�D��K)I�h:�eF|;7s,k�!�j���4{���/�p�{�1�c��S&�}=lN>8��U��K�S�M�a�3Au�:�`�~"
��bB���"�S4M����g�@�Q���im#f.��9m�_�V�;a��<M�ٞc9�+.�91��F�hNO��v-��aXv2��B�x}t�:�*4�$��g�_���E�@/��d��zPj�7��X϶����P@Cs�\��k��#|�-<���Í!�Ecx��5ͨ�Q��>�cW����t�L�ņ���Ka����N��:n��٩~ԟ�ciHȢ&pp��>O@��G�D�ќ'j^�����Ӛ�d��*s'��/6�4 s5��
 ��\z��K�ɂ>{!i��q�d�-j(U��S�G��c3�8~#W޷�Z~�z��_�N��tJ�H ��#dE-R9�s��	�};-�/��K$��1�_�Y�^�_�д��f+����Ȃ��(���s��{#Γ4J���*	FL���TL���o��C��b�?�,�c�F���6-�'��ew�t�S����~s�8Z
�c}�(��-��w�v-#���j�|?��!��=����m���w+q�hx	#��BA��$Xo�~�HH�E��@�O^|_t�P����)����g����v�#�k�ٓ��F��Dp��˥a���Kl��.9��
Z���l���l���Z�)��3�T�DZ,�A���8W.��s�}*������z G��W^K�&�ѝ��5��U({ʽ�tj��:6���%���6r}Q΄�V��]���)O���Ƭ�UO+�E������h����Q�q��|���r�jdvN�,8��H�iŶ�DVf��bco�\c]U�Ic<��LN䀱���t伝��8Ƴ��善�#�Ij:/Yߪ��^,�+	�5���!*a틬7�f�'�yyV�%���J�4��`%��XN�7�d���/SQ�w�fL��-
>�bm
��J�P��gF�-��\b��Xn�����Ee��y7�&���ڂ�a�TI�[�y)`�T�l��{��}�8�����v�]*�~�L�d�}��[�����`��|Q*<�����X�
�N�)m᠛"�y)sF�ȸ`|�˕^V���5�tw�u<:xm��B�O��~�Э}h9�+��*�$�]jՉ�1��Zjw��V�덎yY��ك��}4t�d�="!/���:��q�����gt�rK�f�1Dv�{���6R��*�$
�ه+K�7��
�w�G?)�p�⇈�\��Ԓ3�ꀟռ���Zr⁙D�zs�<|�hH&�|��]b�K�� L���bĨ�͗��u�0%�=�=���#�zCʫ{��c�V��J��.@�d�2�!r����-3�n%�FŬ@UE����^ U�:�A�e:��f�LE�?�>�9f�I6zb�"��w$���x���F9\ ��?�	\ė2�k������0��!�sFO�&����>�輂�J�[;�<��qJ%�As��g5���#�l��s@q��X��Ml�`��By���{:�"�@���O��Y��\=B��_�"� 	��f���z' �]�E3�KGVòEw���)�6h��V}g*{
^@�Y�f/4H��������X��>����k�ʋ��
�LvAq�gHӉG�7�Bg��:��? IR�V3�Iaq�Ƿ��l�@�0�P���sqA^`���h7\ϯ���@���cNȪ���Y��.�R�dsd��T.�����	'�h&�L̃}��n�g�x�N�I�7��v������w�iN�J��C�&$T�b�BS�	'�lv�^�}�`N����ˎ(C^�.���8��ʷO�@�DM�J�Fo��ѳ�rM6��w�$"Nq01�Zg�jl�X2C��Ռ���,z9��vL��n#|D��Z�##���]�Oa�?��~r��bp|2P����j��ݸ:yD[��ͦ���O,$���UI�Y�]c0��"jH��mL��<EĆ��wmwYnld\�q;�����'uu�HG(�-i��/�7+iy������ks�����W��ۘ�����9:z���R��ny�bNY��0��˨� �M��yD��y[v�/��"����%z6�������x3e�Mh2�h��=>��׭7'�X����-��m�/oK�\	}��띹�5�Z�cGP+�럸���(�i���������N��E�Yf����J!x���������[X�V���g��J^!��ɿSU8���[��*4�����Gsow6����R�]�����a�nhǏA
�>�y9�@��Z/X�� ���5a��߸\��=�3�3!� �W�Ӯ�p:[wFٲ��f� �5��kl=
�2QzG�x����B��1���\�8�,ӟ���ޒ�ه���~����3�.[���?
����0�YV����]����9�,I�[*z��kS���bc6Qqh�e���#�����n��:��������)Ҟ󎢺�P^5V�[��r�
f���s���zZ;?��IźM�yM�`�Pl7�S/7B\8��x�[d�E']��p@B�	[�аQq��/R<,�"��;����E�f�tщȪ�c6�[����s���E��Ԩ����S�����U��u���_9s8}�2d(����j��6��g9��/��hDW�X� ��,F(��!
��Mu�-&��l��������8��9�W�^#O�_���aO"�fJ�5%��8�C�X�`�5U�&�
h�b���2��miĜ��e��!q�=Us*۰��|׊�$�xE�GIJ^�O6i��	���Ţ��P=ʻZ0ɿ��(�^kk8%*����Ÿ�8���쌈��i�P�{�
j�l(�IX�MQ�]ف�D�T4t�Z0j���X����"�s�+�K|9f�C���	�?(���;ضvQFo)�u�@*�A��(�ȷF�,n�#���e;뚽��ѯ��KZ�v���	��V6$z�����	$)X^cWh�5E��	�����<��GnϏi��AK(�W5�G�s��CJ@��z�n!:X�N ��,m�3sI0�K4/��"jɴ�uI&��e"I����x���kñ}?]��������%Q� �.����2�TY\�y8h��ղ��;C ��'Ϣ�h��HE��:��sS�#�1�y�^xUV4'��i%��P�S6mj�4�0sP�/X�ZM�Z��>p�0��:7�ڭX�A���}� �
�jO:CV��_a �U��l�}�y ��>��$ �lc�:k�j������`�]"2��e`���YPu���`�������5OV�v��r=v���A��xE �?�\��_c�v�h��Y:��A�R>�������հ�h���Dh8�a%�i��������f�3�z,�D�J�޻Gڎ���@0�N� z鱺��֭�@-B��mZ>z�/x�[�lv��ĲH��v�2m$SS}�{���h�;�,QhJE ˽�o�=�<A�>M��i�J�����[|Iu6���Dc��h����I��%#XE��DS�"h�#�]G
��� �?5�c�N4�4�"p��>26>����0�)q^m[Ύ����5h*��-۪XTA�8�N� ����aï)Zga�E?�����A��b���&��g�'��"�&y��Q�5���4��E�:.�)�E���Oɚٌ�r�Vj�u�*l���l��8D�Z�hi'�%�l��y��M�5!
.����>����4?g���J��=(�z=i��=&?��w�M>}��)�M!TI�U@j(v�\L��<"�$����2��ȗ s����ת���S��.�I�ݠ��3��v�*�@�L�sݡ-м���Tn�섬P���*�.�Z�L�-N^�B�REv�H�Bfq��&ܗ�.�_*�b *}���N�RT��H ޡ�kނZ�wtt���R����� f��@z��R�)��Q�s����P"�ot4_乷�����l���Z[h�В�����f_��'<CUS��@L�B�39jK@mn<�y� �'�F���Pf����ř��֢����3�l���+i�VF*��j�����~ �(�rY�DV���YȚ��CU[5��:��(�+��6��^)�UB�Mq,�8��N�t��.��#u(����A��}a���ao�k��x���������n�Z[�Gw�6�ꤰ��fh���߁-H��~��.\5�hGj"��T����~�ﮇKD*[��"7Ȏ�`�n�W^�=�9�.�'3i�Y�*U�Hi���c������I������"����\�\M��d2e�:{������\;A��S��`�8Rq)zO�3|�^8F�c�y����Eq�i��!.�N}�z���X>&E����UB>^����fb���bS'���:@�+�#�U��i��D�lV�qo��(	rv���Y;T��a\�����ܩ�;�P��,/j?s�W����he�Qŉ8�Tu�6d�s�����/}��H�H�n�D��Ķ�R�@��Q���~�_�t��Q)9�d��dY���y�.Dg����7>�F+�	���GW5����$�o��pȝ՞������1�kaT��cJ�n��D+����M��nܦ_����$���g�*gE_k?t���
⢫K ,�M���~Ӭ-��@j� -��N�묰⁾&�;�+ܜ&��7��U4������m����A����_��u ��b��a0e�Q[����(I�9�	b���IƱ��W/޸�����O��ո~�ɚ�'.s��]2����EZ����$�i��0$�m�����Z�b2�j�X�n�'����՟r�����sP�$���f^Fy���]*����-vP�od����T=����Ɣ��}��v�fEU���?�)8;�E{ϵb���;�q	oq��)����8D�%��Z�6�a'I㑽D���;�;���N2�~bk��G����76�xo�T�3�=#��-�+��s?�u��8*�h#5�gH���=SJ����OD�k5&���)7K1�1��\��nҥ�1�˔����$.8�0BG���U�V(�}t�ye�D�g����j#��9�-�"LY�O$<�����vQ��8S2i��m�Q��ť��
�H�}Q3M
����IUT��?�|��4�9���S"�2Bh8������_��ߡ�[y6��z��}ao)�r�W�H���nPr34/r��8ߗ)�0X��6͛�@
�(193�����V�M�>� s���΋��t}&7X�迌�����DE�Q:��3:6"�1���Ա�}Ytڟ��<����V�G		�$Ҕ@���2�h�u���]o�|PD�;��\�{Y��Ysc�i�G���{@���~��	�'7
�O��b��O���8 W�Hۑ��� �J���Cai� �_֔(�c,�.?�K`����p�u��� C-��ͣEt'sJ�L�:�{�ԗ#FrH��[Њ�1O]"6$�P�)�;�yf�!����'Q��8%�^����P�Fli\M5bVJY��aI�gn�g�<e,!�򠪅х5��s�$:���)�b�"W���h��&)b�,�m'Af� -<���m�!���֬L������=�q��/��cc��� ��3���2��u��S��զq����Pd�~Z��'�<?r�L��u��҉e����e9�	�b���,�#n�����Q5)䓧?���0؏�|��V��43����u�F�:��b�$���dO!�ozIU��Ű��Sq������X��h�*�%ܭ��o�<v5��G���?gg��O��+�v��+����]��,q��T�I�&�j<�ꊫ�9�P�X3f+�-�X��Uqc�s]��H��-x�*w�M:�2�<��ez����?�DG��_J�ްK�~�",�.;�\���H��)��tI󕃋T��d�� `(���"�B�� U���V^��8�0#5��V�z<��Y������v���f��&ג��_�K��T+��{_�J{'o|�i�ӽ3��W�Ĳ_����0��,�3n
_�xH:;l�T3��G�ދ���3���/��LX��o��:5����]���	#��Y�?4�񛮰�ȷ���&g��@�
� K ʡ���-��N��>�f�����8�Dq�ϔ8��G���������䣁̈́�%{GY4_Xo+e̐v� V]��j����=uYj��0���D��>\xG�c歴B�ԵA>'�h��G�c�ӛ`~}��iI`x�}y�#O�Z�^�H�m��S�"r��f����̯��Z�|행�H��0�a���o�
�nʳ�⟢�r��Z5��Z�F�"�k�����+�$D��?	0��x�NŗsQ&F�;}Xp�T �M���9��V��\� ��w`�����:�=`ˏM7W�ɑ#1����av�WS�0/�uF4�p�~|���!my����Qh�c���ZA(��y���TT�M��48<a��dOR|��+��H˚��g�:?�b�E�2�v2O�/8�B�J8�S��<�1I+A9��F�5FX �徉_*�(��]�$	 (����{=KR�/��ʒ�R�Jڞ���b(Rb��7����ZIe	�ޟ�`�G���h}-iӝ[�V�^'K�sߤ��⃚��2�fC���g$��ى
���ⲏ�w�|ѦG�����F��R�\ȴ�@�*�4N��o3�?C���t�&;%�s�D�u�hT/Q���`Љ+�gخҊ�{uI�Y�	�}NV�L
J֐�3ӘY����h�6r�]�����[�����ˁbH�"	j/���M�a�Ge7IK�;-|�Hq�Dډ>�H��e�:�}��� 0���c]lfCd����tz���k�_X�]�^���k%x�!�XNQ[�ލm6)�U�~�Gf�Cu}�jv��ba,�
�4nj�]�ȝD8��2��P_h�=�N�1[ �(ز���R��Ŕ�S�*A��P3�w�o�o��S����AO��霪IO�Hqc!������l��AFy���vi��_�0��d�}@�%X�9)�r���+����M*m$}��d��� ��'��p��\��=gI3vkz��;��+��Úf=��Wj��F���7�2�]���k��^��[F���ӯЬ粞��В��W"H��켕���q=y�2I�kd�>��\�||_e�-���Wt���2�E�Ԗ�V�cO�Y���qJ��̍O��V��� �Q�6%?�E]�߶l���<�D�{\�x��ψ-d���l���cq�w$�e=A��.�j�m���ԗG���ߜ7:�1�����7$~���
��u5��N�(���VF���r�����;W[�ח��[QrrՇw���ިM	ˈ�A�7�Q���h��(x@'*eT:+�V9ϖ�V�.�r���6��PFv���-���.�!���:�%��|��7A5޺Lm��+���)�� �Ў�c�q�m������J�	��L7:io�o��t�~\oN���/w*����\��G�#i�)��鮝R]����^G���;�ձ��+=a3;�����^�9�[����?
�{�=I*eŵ_k-�u�}:�=��(����k��kI
���(�&s��Ԓ��
5�*I��ٽ���Rl���/�j��C�s�=mD��C�����N@���omd��m��qԇ}]�W+��d�0�<�:`X�6��:�d��{�)m��Xs����C��	�Q(��!��8�j�yNG#�������2��ױIW�7.��z��ް�@�n���`$و����k�q�4�1�p9D�8��� ��&n��.�W~�;;�"�=S�?j��}M~�u�|<Cd@KJ�m��Z�+��d�8�BN��H���\	W%�P���.�^~�_���W���#-C&j�sdM�!#�B��y��d�#�ۊ��ǿZ�՜�4&Z=�?���z|%[�"� �<,L#m_�H�|�V��P{AlP�B3���p�N��KR�j��k�5�d��R�a��&�1���G.bn/2�\���mo6�zܮP^jK� �8sF�0梵ӮQuIϓ�;�8��-��>�����\9F�����g�=x�А�"9J�3�Q���7�p����"�=�5��Pa5�ٓX�YCL=���Al�,����H�`�w��Kk�Ӑ�H��X/'՛���G�\�v�%�l�2)���L#�+10�$;�S0���(/(��ߓ�h���D^1��6�PƐ���/���F%������FZ�k��5��Rf�\-���'��F>��i;�6��"T�YP�r7%N(9���â4�����78���g��"���d�+5�x2e�ԵQ��WD}w�:Җ�M� <��)���'$�ɯޥͤ,ӗ&�]��t'4'�qT��O�@��RfC�o�!���۪�e��I���ҟ�����%��G�jFF��r��@:�"����5�>�0�����[b�?��i숱��q pV:L����ͦ�Y�R�~0{t�;��Q��W����ݡ�v�d�@���7Qm}>�1�m���>��ҝ�jg�6�S?��S���y����^13�"��1��S\�S��BKj�����t�B�Rx[�_�6_+�q%O�U���U����Q����󆴔�K�Q�<�:B��ģ0�e*���M��Hd�j�%���u�J1����KM%h{T��P���|�4>����3C#$X�́����1�@UA!2�N�q^,����c>/�����v�����A�� 
�|T���pKθ�5�����))&̺_�4�>N��
��x�`f�(��֦�يb�[1�e1�b+�K?q�
	1���%�D@���.G���
���')U�W.aQ2|h��M��/�"t��Ώd�������6ee�D����=i�<�x�����O�-����(%��]�W�+XE��V�j0���#!���:k�긜�y�����fTdVt~ɫ�%��ɴ�V�FrG��z���`����.�3w��v�ڡ�/vu<�@e���ôΙ�=�K_'[�/�\�.�s*�4�V57e���YG㣌��V E�so���DJpNz�HA���[�-@��E �n��Ap�jhcp�uF���|Ibh@~�K�i��M�y�e#��wKػm���N��{V=+��b�kJw��j��{����EB6�%������ࡻ��]pZ� ;]͵�*,ݓ"$��ͅ�5�i;��*\��99���>�;Y��z�a=�K��+ñzծH��菧��X��L���\�K��Ǐa�h}B���F�̱&o`I𖶂ɮ&�6����*��E&s_2���{xt?�vG����ocØ��fŌ�4:��/jQ�1
�I�.�~fX���M���;.v�X���D������L�
b>� �/�00(�ڤ����Z�-���z��N�iaNe;-�"�7�#��|�Ҿ�L4 
:��hC��X>F� �j2��NP5Z~�ҕ�R�������ۻ2�n��8SA������L�3�.Aܖ���m��q��v{����}W�ç�I�$�q}���6�Y�P"ͥ>>��"q��"@Ú���9��Z��d�����	��І��wx�o	��O�ethqr�c}�A࣡���Fu�`A(B;}Pi-���n�xd�|�v�^�ǬL��R�ۓp��pV6h ';�>��M��~#�Hހ͌Z�!:�h�!�:�naY@^��[T��m=��U
]}�x��H��*�|�R/Ҍ������K�{��o2�u8�
_�����9�wW��刽,��N���r�
�ژ�u���T�=�*a%��"�@��qX���� `�A�d�7h S ��e�Y��լ�2����\�����Aㅳ��0�nTN�����̺��e�(
4�B����v� z���G&�嶡n�(��+� iEK���.ߊW2q9�[m�A����Mvx�����{h|��e��|�b%��H��h�e���H��/A���o<�����knݫ�O�ŕ�|�
�RN��A��Y��Z��留��KZ����4�|U�%����|���ȕn�Xw)�G�ⰶ��V[���h����5ge33�B89�s��[��&�9=�ҒI��*��]�)���4�b��I�]���W����z+ r�ї���F)�⹕�VRf����%/�]���R�fzv���~
�ȏ��C�J��.��l�5Ć��{��U���頫�|x�_�'@�1襰�QЌ�~7-Z<�ʯ|w�!����U�4�qzﳟ�=�ثW���؏��C�:#� ;�]~m����T7�R���D��rV�HK�8I�b�ኊv�l3�#��8���u��ϋjɪ��9��RhIk�~��9oG9�RGt��f9�����ė�E�<(�Vxø�����"��Kk�|�D��Q�Na�(�Į�k�n+KKYH�#ޭM��bX����*�f����,{��8Q�I�H>P�����z�F�����r�`\ 2�ۆA*8�&��L�~��&�̢�����7@k����͗{��߮7�{G���w�O�/}+��Ȟ刧��,q)����X�������1b$�f�د�ש��%�4S�Xj�&�\r��/,�w�A.����v����_��3�ȏ<CelI(�>��M�F �DHB'4��ɖ���C��x1���9r��4@F.�8���)��/�V������?��0h����)Q+��egَHDU$ϖF�z�M��GV���W��_�k�x��B�ES=/�FC�N�d"��:��#ܒ��(���K��v����+�_x��m���C^uo�{p����8���ߏ���K��)�Ki	�i����=�2�(�c�w�߳DOL�� �E@���ڹ0󼃆� ��,8 ~�JZ/p�O&�Z��h�fr�R���z&� G�	�膊��T��&�v	f�=��;����0xω�5�a{�p������3_�k����c��+`�g'7t�)'L�pW���Dh�O�[�>v�z�#턃o��&�}>���7D�!�%j�N7_�#�ۨn��׺��Y��>N*$X��0����T�H��μ*�� n8�<4����m���n�S���D��@31	Gt�LZcj�z�uW	���Z-�� !��Z�E�Ń��~p��#��.dMX{d<q���ho�j���zq)<hZ�%��KF�KƾV�%��v,�.��y�F�m��N6b��i�a�|u�2, R<ZS�v�r!�
�����N��&����v��n�i��ʪ��&%������F�y0���}��XHo�C�D��㦥H[��ʓ?�^�h��.�|1tKm���E��Ð5���~����[�HCd2���>mE��Y�(��\�mY�f�r�zWC��e�i����)����i�2��xTa�`�����8H�R�pF�f:����-2�@�^���*o�6�f;�$��k�q�ѐk�qp�~g^����Y6���@q:�TV��"�$_he�3�c%����Pq��^Lںk�1�T��opI-�K�V=����ic���6�]�Ao}����U��YǎR"�ܝܕd��(^���Vpp������)e�ڀ)�ds�GX���$���n��u�J��Q��&{��T����R�e^�e�9cS4��ũ�mb{� o�I�����U
{&<��D*Ğ)�;M��G���%��;+�$;mx��[i?�瘨��e�4�3l:�`S��"�˶��/����p1Dz)�_�_7�F����h򛢭��7�+��v��e��ϋ}��X�3�����s~���_U�K�l��p�ûlC[�Hv��,ê�Zʞ���#B��h~�,�W�p7^�T��0�5���A$#9��=g�B�k�'sY���L,	���Z���F�&��lp�]��z���P���[q�F�N���w��E辉��7����3_�a^h�j7
���օd	KZ��K�A��[9�i%��U�O�<�w]�.r��6�eQN`ɵ1B'Ȁ3?�9:�2��kоrSŦ2������W98���@�����Y!�/▂�Mr/���Y���%�)�n�p�Ԡi��%r�Eh��e�s�U'�?�����^����_�A:CC"�^'����3&��Pjz�K[:�)��������+A���{��ܣe"��᭍���Vg ߪK�M���<]���	��tO�*�g���(�����v3#'�j{I@@�X"Q9n�#�#�$(����^����4Р|f�Bg�������vk��V��#O5N��?(�%c<���|2�5�n
�t�Iݸ�X��g�`���ka���Xw#�0���1����%�*ED�nS�%��p�M��`u��4���Nge�h�L����&�:F���:uT�LxކcjYq�^����Sl��ԡ[��.�|.�tr���je}���xg(��xDй+�j���7ʸDX���Q�(�D܃o_�.�G���M4���?1�!@i#0��y5�pA�%\�,�ƛ
���`To����7�[� ��?T�Y���ˠ����m���m��w~�~�Ύj^�z�(���Gy�}��"�Ͱl4Bˢ��<�Đ(�~�"�0�)�k�c�!Yr欟�t��hu~�P�my3��_�:(b�_�����t�R
���RH��w��A�7c�c���3"��+�'�HI�򛒌	�gZf�</4�HQ�-��M�lj1,9P� �!��c�j��Jc����;�2�_��Qf��S�ĊY.e0�Z��k:b�1k��$%���᜷��\IZ�ܬw�goP��f9I�V\qH�	Ͳg\��U����`*��2�ۨk���y���;�I�O�Ѯ"W	�\���r}�2���#�}4�4�"���3�j�BHΖ�u�APF]�x
��`����X�8.ج���<����]���fL�|Z{��3�Z���2w��v���	>F*<,e��%�}|�J����dїu?e����&�Uj�
���Y����A��vV�2E4[A{�Z������������m@�?Y<�p�+m��8�Ht\�	أ$�O�?F�Cm>�nũ:���{r�ܵ�g�ǟ�ߑm��xE�o&�/���p��}�$
�;���T�;J�2�8���_�K�Ͼ�k�\$tO(�������d΋�� 2��)h�10�W[>L�u���++���ı`� �t��j(Fj�3�����D��>r�H��נ@��oX�Xn:w�]#R@��d�1"P�;�mY���%��\��Ժ���o�D�3$p�ǜ|��3��k�v>��'��S�rB$CDE?���7D A(-A(x��G�t�5��}�A�^-K�P��XVvz_�[)�%i��edT��w����4��ϒ�ې���Dv��.�EQ�	D�l���}��!ˏ��'T�P�����aw'�����	W-!;�}r�UF��\hzs�$���ԛ�b�����S��
�pS��Cfd	������R��r����	��/]���(T�s׀?#���G"BSe�7����3�dB�Ô�!�2o���0?.�v�Ɲ����+}�S愆�y2�s��R����H��l�+�q����Y3n��4l�%���j�ˏ�N�V�Ñ�ؖ�$z���P�**,M�q$-���f2?�nX�q���۴��բL���n��:ȇ����\��,�b��J�W)�
��`��I�y@A��� Ѐ�
`��]����gք�Q��L?C��
� ��L��Ġ��C1��I��6z��J{ܙ�I���e��f���E�VF-���w�v��6\�W&S2���-1�@��# �����M��Źx/�H���t�^]�p/�L_ַ�W�k���NUqs���J���,]�׸���V���zr��#��+�hr��9^'�X�nMB>ׁ� X�}V�:�n��tXb�f�����M����47N� �q!�}��M�2y!M��=�c�"�cT��J���h����Y=���$W�m(t
YR��ߣڻ����)�l�-к1?3�������*d6{"}�#�캇�ġ'��x�-2��)��{�0��fcR�IL�,�Ө\]�X�mhI���=4��m���c���;|{c���\���"�9R�8�~3��J����z�b4#�����Z��]KuZڟ�O&XVt)9j�X��f����0(��#���s��p��A\�M���,���e$�NM�.�oc֑砅+O���/Q�lѱ'�:�F	�z�g@n5�E��acO�fOᾚM���K�$��ӁAx�ޔ��P��I�9���혮�ۙ�bk���2ܪ%)����cƞF�؁�W]&�U��I�KT죚A������'i��p8�)ì�ĆW�d��.��ҭB��U >2����?G#��ٽ(,�8��P�q\� � ����۳� �����f�IP^ߟ�q�T{�d������X~e�Z�i�A�U�0|1�z�8�����)���Ӂx@$��T�s��a��2^�wQ�z�޻���cx�,�>�NXp��W��}������ة��'��9�`��]�m��W��	�_��~8w����l�e�~w�C�Q䏍C �b�Ol+y���"v������x����_[�IMc���j��vM=��qU0o��U�jH��i�[n��I�T50�f��9[��n��<9?����a�b���~{0����x�V���p�gӍ\JƷD��"��i�����C6#�材�6j"#�!ۖDJ˖��p��#q��Q���)����N'<��U;Kʣ{�����GfS�Rl�1m������@|�����Yzy�hQ�ᢤ[;Fݭ �:�Ƣ�w),D�L�v.Je#	�b�<A�Ȩ�]��,p����"��XЕ����v\����E� �D6js���5���~�]�3��i�
Vu�'ow�ض�-vVt�
V���g���䖳3wҵ�s.ʢȠS�%�lU9	�b�
JDNdJL	p"P�����i8R�F��'8В�[��O��jP���-�����ξ�6��W6q]� �:����n�L�O�p��Y���[2+$ j,�(�k����Eo9Ao+:�Y�(ا�k��MDp~�� O���t�Cb"+�������ߤ �y�=��p��\
v���5�@O��K��:@��W�knp� �i8�� k�٤SETC(�O^��խ����
m=���G1u9֧L�j��o�C���Kp���PO�b�����5�UyЫ�h�1��o�6�CI�w���EE�?g���S=�6e����
��&M��u��-����2|k��s�t
�FNF��;���K߿�����^S!�=��������}"�=�4��F�����F~�T�Tb��HT�,j�"�^1P�NzTf�u��"sǷ�'��"hK>�͘+'�XNa��ݮ���$ �<� 5u@BV�g�cgv"���eb�Z֩ڄ���pU�s��kz]�i$��[Tzu��j���_e	-�8�w���!�>v޹�m�)`d���^~Gr�5�Dr�G��.eb������o�Vzxj�8���m����0��Dۀ���3���hB�6OG�2�wW�0�P�W�B�c=�0���<��!��{JDyS��m��ݎ�pټ�DM坋Of�ye{ϋ*K{x���2����RZq��^ߴb�H�a7�T4$R�+�����-�����\�p�5�.�+W ���Y;;7n�t �����U�������zp��L��0�m��~� ΰ�vB���Ti_u6�N4��;�������Bb �����@�ڒ|?�P�mn�~��Nnn��ߒ0�Y����bD��yO�Y�t��\\LeƩ�-߳�b��iAE��s1�٬d^(�^��^��6Oܱ�CٓL�\)�c
�"���3 D��Q7�Q���U9�a!�-](k��t�!e�֓x3e�ަk�wc�]���G�(QOukJ'B�/�e�yl��)�]����m	��_mr�l���f[z�T��n�jd9�y�`��ɖJ
���g���'0�p���<�����&}X&:����0�9;5E��Cz��#����C��H���U���-'!��lļڑ'ɕ��A�o��w����␇����c9��[���Ů��J���<��躮[Л���		r���2���U�l�#K��)�B�j(N���+,'�P��}F��g�\�x��fzFiM�
1kJ��� ��h>_����w���
�� �f�G�l�W� 	��4_P�`�oNYn/����U��6O^���]p��/�"�G���1��(Ao�zГCSI7~욝<�Z���K�#!Q��6��7g��ƥ ��
���b��)�{H���pӎ��!+�TX�1���[%�����50�ԴTT�!}�z��
��󙖝s2ps`��Tp�x6,t\�ld*�bc�����0v�嗓���dB��R����'�<B��:[D��������0��t����Q�/���~�d����Ā�M�L,�6�ؗ����r��v�F;��Up?5��Z�����wlT䙞��G#�R�TRY��B��:M^�ƅ.о�Fw�y�x1��qc=^�aI��N��GB��iXH��	��d������# /J'`����*��>o���$��mvJ�U}�����n�����˅
��
��!�Q���i9v���p6T���L�X3z�� PE>~l�N�N85�PcL�N���ˏ�S�\�du�Р�E�SP�G�lXӘ�6��h� E�e��;f��]!��P���o�<���`����Six�
�ӽ>��0���r�u�L�
;��'�����;���f�һEFO`��o��$dHT4����܂_�_em�3=v63��a�hE^%@0�B��TɌ�v�a�g Ĵ���ѷg	^=�u�qP?}�3<��G�(�|�q8ֽ�תY]VQ��r�u�'��@N�|lY�Er���u��}<���"{�p��+�r�=G%�\K׹9+;���I;=ō�*iI!��R|�B$ַ�[安�5�J{R�1a=�m_���k��Np��7��X�#�����æ�����Zx ͰξFo���%����I�N��A�Aw�DGA�-\B��w��j��X)����aї	P%H�����v��[�O��+/p���!%j�Ġ!����7w�_�j&��ƄC��@j΄��T��u�Umn�� �_8��f��-�|�Xl�A��L�ЖI|��XF0<�Ɉ�F�YS�����|F�=G)0�Ւ}bG�jզa�h�.�F��=O7�P0({�;������<W�_ݤ�Bk�$2葚��	�fU�������W�D�D�Ptg��>+�B���/�d������V�Ů�\�5�-�����u��N+~�J	��Q���b+���e��x�O��6\
��4:��ډ�،�oyq/ƅvJ�\�y��(:Y5�G���
�����)`�Ki�?/�i<�c�ѝ��̰5
zwH��q�$A���L7���ׇ�>�������I��H,�i��<Zi��77b�t����G��l�&cY��9�%T��^8�B��J����Y�<B��T#냬�۪3g�%ChxF�� E�����{��"�	�4d�/����?�P��K��j�Gq$����aJ�8^��`"�!�������J^Oۜ��cm��HY����BAa��i�ls6Y��ڍ��0���l�|�j?~��;��M��-F
,R�����c�;Wai� ���������R֑���Jz݄��� ng�^{se���.L�O��`uV�nU�*}�a�	���{�ݶ����J{��I"�`г�'i� ˠ�h�n����K�ܛoCm*��±嚂o6z$E�
OGq+����|��ՠ��vi���@JɔY�KW^�C���M��-ld�|h�#;Rh]`��u�X%�x��$ҔcJ9hz��D�����E��V�vt&���7P>)2|�)�� ^m�E�]�͓y�䧗�A �(�ÀD )ѿ}dݣ3i .��|w%|�e�2ǚ��tw�����;��5�R��Jr��r4[N��=�˼��-�$�����h=8�9��J�����W����̿��$��P(�ĴbÆ�-�$l�8�Ω���|����i*`��N�E�F�g=��'�D݄9U��N�D�|<��%���mY��)<��g�ws_�ZW�S�>Z(�^�;0U�@^��J���H�t�.?ޯ\�KD!�����oJЍ�A5z�*L�iǣڙ?T��'d�u�u����!	�}�-{T�km�td��ɫ�a���V��`ԓ���-�p�V����w�a��m����� ;��LDK�L�T�6o�4��������Ձ'/J7�`3;�I��4�. ��}g�\�r����nm߬3�q�g�O�����C,O __!���S��u��F+����Ձ�Rp�`S2����*�����q���Ti��{�ur�Vv���Y���2ީߓb;끡MN�}�Rj���=�Uk�c����]!�B� �V�˅Ɍ��U����e)V�6��[��
i�&�̷s
��؛:�&#ek�fyv�Kvl�5	�oo9wx�C��ˣ��E���_B�<��]�c��X��f��r'��q�M��S~�^�?2����J��3-��)j:J�q�aEH��	�GI`&(�o� �r��P6���G
�'�.�^o���&���6�Ԟ�</[��C+F�$Bs�]����"��mU�ƹDl����r��M|�<Ѭư+Ѷ���i@�lwGR�x��$Da��'�u�awB���#�j�>�Y���o����ɓ�x�Jސ�Mx���ʾ��X�F��D^řA~(�$�����ܐF�o_�RXg-�-^F4�2
���"I�-x������Q�s6����2���]��o�Ln�~Z���o���6�`��^��a	us� �2���gyk�_%Q��-���n�i�h��z&kc]ڄ���[E�;!�X�"v��|�ul4<�/���]�eZL�)�1��R�ލ���q4F�4�G�PP�[::�2��,YMs��S}~��4�P	\t�d
��ZN���ω��w&��aB"�~G5a�4Oţ;9���?�Bg�[�fUFָ
j��ؿ��C|g���^������Y�Þn^y�I1	FK8�!�Ɍ�X߶��JǗ2��_;vŃjnȖ��
:"Hv������hF����L�{�u��!K�,��~頻�eZk�+HYNo��kaQ��f2Z�!�Ğ]$�vS���$��L��ɗ���5&�U�:�t����P>����y�*(%|�f�aimg�vn�����`C��6���W~�a�L[z�H�y$��}������.�w��v�G<��T)s?�,K�I�33ؗe�\;�Zբ�g�	�"n��i�'�Rfa���`��!���A5��]��G?+F��z�~ڍ���y��be|j���uQey7 ��bZ��p����(q������uP���CjJ1.���L*h(�*�J�Q���,O�����3�v�+c(��5ކ@U��%Ҩm�&�pjy�Q�
��&`(�C'�?�{Wc��T5V��E���<��F��X �m��6�)����0����)�7l j��܇�ǸT��c�Z!��B�x�;�5�G���^8��I�A|�?��6�I�_�@������?<���I�˗d�05��/���ӧ�@�tGYP ��;N8��~�ZqY���u4��(��R�B��*"i�Zߢˀ)�t�}	���b��e�bx�w����R��W�=�2���]��
�,�=����������Y��E��	�TG�E9�_wX�o��d|PO�=���db��7V`4�'��Շ������w#s���D��/�%�rgG���No:tP�����i�3���_��f�iW�|WWH0���Fo�����#f��{��F�p�iUP��2n�}�Tk$j]���S�Jft4�&����~5��VI}k{K�@��%���/�~���~�?��<>'�|�s��*lzV��bJq��Zj�,*�s���T�Fk^9��B!!3D�����n������@�$Y�Ξ�Q]��򌚨��C�e0V��[q�T ������FB����6�9�C������h[§�^�e��t�YA��<W^J����+8(���xOp������m�?�{V�$(��C���[����X�!�H��[5�������%�6#N��0�囌 Rb�
ڻ�vߤ�P��z������0\�Զ�}��+�je���*h�Vt2r�\��h�\��$3f�^hQ��&�.�{�N�Zta{��l�/]B8�U������1$�����ë��Z!!�'��K8��V���`�M�h_���_�rw	�Q8��� 0��G4|���f@���v��r^�>X0T���0��Sx�|����6NJa.9z>L�8�X�K���3��Ck9����<ώh�a��H�0j�rݘ~{�g�+���d�g�R�fWG��@�傯��\�y���?Wmw����/�R�i���sV��#u��e��U{<��n�X���T)��9���@�:�l4�{�{[�Xؕ�$�Fдp�ہ�d���9i6�G��;�ڹYj��;w�z�r@aT�g�Y
B>E4����!��'A	�(��=B�4����&�G���T@8P_^��I���@���(��r��z"�v����73�Z沨�
s/��(�`�'t��_=���u���W�AA��	�w�=r��ө�P����ɛ��>6ʁz�/���`�����*�1�ٴ߱���"��l�y�
�ȝ��� /~�eY�MԦ��֣�xy��H�	8T�}~��O�a���#�eRvʷS���l�a9XhԞci�+ϕ�[�MD~�Emr��m@�ևt2?T��t�䉥0�֧�KC�������
N�H���*�;wV�.^]}R�g�����YM�?���&ԏ ɮ����W�f���1g��ƭo[C~�0���oRTFK� } �y�~)����El]���Mx�*���x�@�ߗ0��s�&^U�?���҇p,�wW"���)��3��W8��l%�w�����N)W~���2�6�n��$'��������Շ��VN�r�#VM7)	`ߣ��5�>?Y�A�$�G��2�t���Y�����qE�ZQ#Co�1{/�Ǔ`iw]zA�
����<!�:�-페}������te9��VY��%�#�~��ᦳ���o���@l�5�'������ ����S�˂��g^Z�j��C�׾n �Ii��R�|#�-9�89��Fd�mQ�ЩI�{Q���1��خ�>0�P;���C�",��Ǹvf�$�6�f�U9��쁃�S'SQ�\�G	_�� �wob̨� ����	N��U�S�W�����6y5�Í�и,���� O ț�-�C֑' �Zi��A�2_^vǈ f�&�*X�Y�%fC'�j6yd�9�2����\��WT��@��#���^D��	����뼼��a�س>
�:�{AZ҅��i^���]��(�o�/��96��1�j���zETˆ��5wO�j�Ə�䛁����aw�^s�A+aÚ�sSG.�������m��z��J���1��+Qۻ^x���L�p8��I#r�g�Y!�$��mT�u?�S�m4Nz��p4x��6�F@��h�x��R ��I�<6 JsPn�T���3���"�B� -����C����+^��H��{�?1}N\øCy��톘`�-ӭ{Q�p �>�WL�'��(U@�g��T�ca�$~ffM.�.�S�D%GX�i8��!2Թu�����A�}pt��R#;��ٍ�;dp���1�Х��g��@Tk=Ȋ0�ˢ�_�9���
�'>t��`#X�"4D_&�MEC�"�QR�*2�Nn�����xJ����E�tݢH��ڪ�� ��軶���Pi�����]\c�l�y�^Z���
�(=����/\Dn���>s��V~�-h�`�e�����iW�8�W�jW}j^6,��T�q���r�3��YlO�aZ�aMZ�$�>U��o���K���e�����w__�i.�?��+e�Т�-*�܂6�O��_Q��^~�?L8u�f��=0�nV�I㧆;-��ê��6�㗰�<+�}*����P�Oʇ���=?��yq~�O�?�0<�{�,���o*�`7 ހ�h�ؑ�*!y -Y����)j(��!��Y�݁�n�t����w��d�hS2����A��mXݢ ��[���鹟0�"�p���Å��z��zk��/���(�gզ����7����tA%�%�9
3U�_|Vf2+֑�,&`z���WZ@���r��:�[��x:��������	�ő�ܟSl+���uU�~\����{��Rq�rz.
eǩM�,��5)r�����'�GOw�y|v2!�����Q�|�?8���	�S�C�WA-�1+�Pz pl��d
U@R��:%�����mE��WɝUf�zGۊ꼙�]*�A��WB˩���J����8�U'��\��W��"V&�p|�I�O�Z�]��� �o��6­����|���a��BD�B�f�,��fB���M�z��A��܈��PaR� �@?%))R��p�+�����n"C
��&~#�	?�����I�o�Q �n���>�h�{f��I��\4��'h(�����F�6�Ѿg,S#��L�T	�=4s���O��v͈;��[H��C�����@��(B.�T��a��g9f�!^I�&�d��܀mӑ8�8)PO�����p.���'V�RdF�}�!�ؗ,4�?��)!���w1�x��(UýB>��B�4���o���n	Ʋϔ� Y�����0^�k|��/��nh��Q�`��ԲV
�����2��D|(���ihG;��E������S!uy����'�?W��b��L��d��ku!�6:���-�0�P/�W�$lu��p���^�ȿM_�����>=!ƞ�����H�es
���0q�&�ȿ��{�Al�;V��B�����nv��8�k�4��]Z�2��iM�3h2M�����bS�򑋴��6q鞦�տpnY�_�
����~&���o�cӑ�����w���&�찱
�8��x��O��§��ߢu�>s[�Ǔ;���y��uh�(� �m/�#�E�R?�|ׁi��=�圀#B.�������Ĕ�h�Q��ı�e�	c��ҵ0N���-�g�G!�& @���˻UQ��1��ţ�U*�+�>T�TF���NV`���y�=~r-?��k� Xy�9sZ��F��P���U�Wΰ/���aZ�*�߉���{����y�_������RQGW,&���"�cpV��-j�	���/�e��t?�V���7��|��Iϒ���m��s�rs[HRhmj۽��e�h��Hn����{N+���b��~F���r[��!g���4�� �Q"F�{����@߻��*�s|���W��L�d�|Í��њVPdql9d	)|�vQ�mķ0��{'�R��Iu=#��'���cȠv z�!4�����W>c�bs�O���Vc�l�E���� Қ�ǳ4�l� +	ꊇS�N�[.j���nw���GH, <z7'��xi����I��y�
�ל�edS-��@�6ό�'y�5�>�'����0F	���/�,��`S]���`xi�b��s����R�Z����%N�H��Z�1�Τ����_�N~MI8�X�7H�:�)w�zAY'��f�YY��-�F'@t���SB��W;��\f�ul��|�`-c���yh=��N���uֶ�1�]鄘i;�F�Ff��v��B��ର�p!��Kzd��~C�@l.W�MWY���t�>z5V1�^��y��(�U�f�<�y����Ծ7Iѐ�>��a��?ۚ�蚦�H���t�� �)��G��f���ޙ���zm4��O����z�@6�ar�@3~�� O�Z�2%�*����Q�ۃ��k�b�x!Ə�c��CТ���՛��CMۂ��0՛,+x�k	u��� �Ɵ��RU�FQ$G@s �,3x�E2�R���8�#�QDM(���H 8>�E�>B��4�>�^.7�"Xk$�R-��)'�ܿ���l��H��|k����\�4wg��B��Y|�}��XrA-�n�?�?�R��BNv���$Z2!~[@x��?r��g������5���S���Qp��xy��T����kS���ǣ�p]�s�Q������lE�J�֫0Av`�>�°� ��"܇rJ�K9pfܽ���L����*��UZ���	7H�aI�`�W�Wm�$�_�W䷟�*�䊡�W��v��M���S�fF�b7��Qp�0���0`n���>�ڒRy��d��in夳�>9p�bB�ֻ��H��J������@t������G����c��������m�IG��'�Q_��!7�$���~1vo�OVpK4���:<��F��a�$��h�D�U��w:v4]����/J2-@�;O��#�e]��uF�*�W[����'UҜ'�.��2I7�Y���F�ir�*�B�v'�Y�����/�7A��<�^U�,L�;��Y�	C��k̈́����S!2+y�L�Q�Ǣe��,��>�C�[* "V=E�L�;k� g����@��s�� �*�����+�*��*P���13���X�J�x���:u%�#5���ݯ 	M8ʑ5���X>��J���&�dA4}�)ŞTM�-§d7��͒J��\�F�DC��o���x.�I��1a{Nmڏȸ+D�J��������A���5aP�eb��2N���\���T�h�ˊgŁ#���zA�(k���ΡJ���<��Mw���g�q��`�9��g�-Ť�׊D�[���Iel ~L����#�dw`�Zr���F��Þ�����D�	�V:{�O��Tٖ��c�s�-W&��$) ��
�GȞ�]��O/��*�&��%_Q��,9b��Z����^U�:�h�P(Dn�Z��	/!\ �~�wm>��`
|�Ko�/���Xոp�]��g�������/����f��\Z�+�FD���vL9e	~���B�Y��.���m[���� A�=V���l���Tm㊓���G�迵u)��,�\���U�8u������|��\	yJ�-+��p7%�$NG:u����4(��rt3����W�)�~���E)�Y�ިh��SO���$����7�����Kk�d��KK{0]�\�F���be�~����c��ۛ���|L#:$�q�+qB�zj-�-Z&�J�X㸵$�{�b@���i�2�ш�H�>'��
+o./���_���nXF�b<%G�N��ɽK��0R��D�ҍ?�!�&r �t+��# ܩvM�oyS�j]WW�W���r��7�q*P�ڟ�J^x�h���ːlOiP����&���P|� �u���h����#��C��i�%-����QE�}�����]������ԩ<��1�-f�|E���Aglj"���|^9ĩ���|JK��$P�@��h˅�q,�
/��$L(%�p�!�d�Rw4w���h�)�i ֒9j@3p�jۻd�G�r��9�H2��|_۔H0��������M����$^d�'9����6i�]!���67�b{u�����dd��&�CD.~�<d�|�+1���耊(6�>DQخ���L'1��Q�=�6%�+����-|�n�8ހt�K���{�ٜ�2 I��0u@�ѝ.��"���v5S6�UᅹI ɮ�մ�(E�O-��ɞ��C6j�沏~��̵߈���M$fQM�6���6���`���7����㝍��Ʃ{��Ot)���xwl�qZ.OV���6���&;�(��+-�v__5��j�œڰ�Q���c��<d]u�}9!��G�3��6G3�Q>J����!�2O�vz4� �o���-�L�Ŏ9�qQ��:i�b��>N���"X�⎂t��Y�7���rI^Hjh��z�
I�oS�a�C��8��P%�ѹ�dvP���I���)l~�'����I��
,{�!k��Vxy�����q^t��6)Ԕ{�ks3�"��+k����Q�ӷ����O����hM�;��B�����Ѩ��o�°s�@T? 6�؟CZ�/YL,`3"˦V�	��t��΁�F����o�BĔ�V ���"��哓�B��8'2��f���$�����҃�{�����#*�}}i8��Ȼ�H��*��C�� X��x��꒦�SN��x���8A�1�:\�2�s�I�%#6��5U1JP�{�����r����u  �=�
�~���@K})_��bl��q�w���_oZ_�&dR�ϼ��T�'q�K��)x+x�b���.�{>�yԘ��� ȗ�Y�$�-��yj�����$٧�Kj������ލ���˶��m��&�&��0)�R��
˂%�V���E��P٢
�?rnc,�2���Q���:�ޕv:�R�5���5�������/�}^���~Ʃ��F78!��{cz[�ϒ�9 �~�#�0U��Ss�_�=3���!Y����0���N�Pb�����V�8�vX�
2�7#^���0��#&V��� �����s�A��{�@Q�OZj���yT=I���0�gi%�?O��������W����M<��@+�&*��ѿl��76E��e��� �FL��L�{�a��Yr��+�_F�ջ�=����[ȿWP��<��D��ԌS̔˪�ԋ��X��,^��	CqZTa^d��xغ���E�n
l�)��u3#U��{ְC]��	W�!`�J���i\�r����<�f{�/7���t�����ؚXE_�QjU�
��ʁ)��]c�k�XS�<���:m��\���T��29��5�mP�-�S\h��O�%�W�A��P���+fmڧ�Й�ڀ�̍�5�.Qj8	7��)׏�$���KÜ��c\��Ѡ���Ү&�Y����0��Z2E� l��R�hD ذ�X~�DN�um J>��W؂v��k.va����Q�K�v̣K�3���$��9{���J޳y��C��b�!m61{[{���Z>���=��nVkKW�Vqj���r�-�.�Kw=D_�F`>MY�|�D��9�,���i�8y6(�#hӨ'�ܷ�9��2�&bw��B<�b��y�������*XfNcTF�9�G�Hwwe�
j���t���Wuܖc-N֓L�_��	o�p:�C��7���v�E��}�Q�?��Z�zk�{!�#�It��mZ��3Q�	0뱡�mL��������� �1U�	J��@c�����	 �ŗ��U-��:�5���Ru6�T��	<e��P�N_ ��W6��j���U�I_�]��-a��d�����n6�16�U\dƀ��zx�ƚZp܀�%.�,-��X�f.��")@�AF�A�Di+��V��ƶ5����п��M6�΋*���k4��K:�8� ���D�˥I�Y .�/��@<��<}�I^������/&��U��{I�褯��3Կ|Bv-�cY��Oe]��K��sP�xW4=1%9.�{�3�J,�m�JO<������=�x_� *W��۰��z����Z:nM-��Lcצ���n���Xͼ��$u�{"������ɓ��>�S�b8�Ϡ��|��8	�FJ�i唂�2�"�����;��+��|����r�;���>l�x��[Ҕ�;,��C�o:)�~ř�%���_G�Q\F�}[x�PN`e�*���ϩ�r��ybj��;�����&ʈ�z�6�����$,Ki+r)�̄dc�h]��k}�yI��9)������DDd̨�w�>�2@&���Ҡ��U��יc�kmiv��f���+�yz���c���y�n��ZFGZ�8���*�B�*=KEJ�G@���F S@���T�� Z�8�?�ָ�Oi�>8_��s�#9Ѣ��|�"�~�!��iU��K�m�s�(]����h6KQq����E�'lcEC[E+0^3�U����	�DN�Kƍn/[�F��<@���|�h��D����J]h�H0�����n�iƃݧ�y�d�(8�� 
![�"�s���&�!�0P��Q�JA���`�˟]��o��ċͿi�*Z���O�X�/ȏ��A�c���b��Sj���C�۸`p��7Y>��1{>V�ˬ���&e/dY��%9�����zc�|n�xdẉ�����9s1�O��Db�u���Z��-�3ɠ�I��Rx�Ʌ���X����K��Ir�s9��)�����Q\ac���{1�O�40{I�%N Sc�P>��L�A+(8�<��oK�;7���೜ @��D�hEm���i��){��4iʘ�=O������D;�*����Fc�l>$�^�:��(��uJ�l_�g�i�	��n��v}2�>k�iTG	���97�mzV�Yj�k�w("Ha�ʎQ�#�i<��s�ޫ@�[ӛ�)Eo╰��eCǙ|�6����y�C4Sa�H�J��f'	�ˮj��{3�c+�a*8�I�_���j��T��d�^�?���A/���\XL������16T�1����HM2��F�E�k5ʂ�af�>��P��U�6{���0�_AP�~���ab=	�]O`�����	�ba��~-���6E� Z[H� ��g�V'��0TEZ�
��]�U��e���?��z:7h
�ׂ��l3 Ğ`9��u�u}+��S+�aF�b>'A�+��7m���[��C;M�+��Lbjpl)ç��,ji�|��pO$������-!'��0�<>#� ΢^�]�>��n?'���q[~�%�u�65Rg!&(�T�E��S�5pU�m6�K�%p{CB�m�D��d��h�	��RF3�危��~hn��<�$:J,�^��,ҿ��ՙL �&f��S �E,rK%[��$:���B]'q�D�0=P�\�]�xnZ�R�6�2"�zШ'9ι>���c戺ǩ��]Ć�5�d���I��l���uu1l��?r�c%c��V�zH�,ɚ^#�o�,�������I�y� E��b�N�󦝿λ=ho�O�����K�r��y���1!�[2�KHp�!D���GX\[�iq�U&5�?�	[�Jo*�7������m��orz�8~⌓r��*����'iʂ;�X��YӕM^4G��X���N>�*�rځp-��+�΅b�뜨fE���<볖��Lڤv�ҡgp+Vޭ��m
%�k��$\��)�X�!ʤy�i�p�)(��Y��ՙ���_�֨����PJ��f��w�"���BD�"]��lNCi��۩V!C�;a2�s�*CLN�"̯	�{���-!;���La��0��3�~�v��S����q��RM��uJ���'�Pd�m�Y'ќ��,C�E��	G�M��G#$-	�<5h�UU9�������D�Ѣ��D�^���g[Aq	�g/'����o[���g0&7���oYkW��K���x`�o��0��<�Į���_�}��L��7������y���I�}�6�Fܗ/!���7_^?�֯�F��%C�����a�S��6Qab����h�[(��V��D����?~yR�k%���40����y ����6��B�Մa��m]�&)�v�P��|p��I���"j��7m8k�P��[w�#x>�6*�Щ@�MuI� ��Rl�m;��7�m��@7/t�\��40>��(?w�z��!FT����L�5�I�9�@��8��'�{����x���:�D��3I��T�ϳ�ވg��M�o�e�� �$a��Lw


��X�x�����I��h�E��a��hf���4N}�V��;�	_9��(�:(��ar�gX��8��=�+�,Z���w(�U""����[tÔRGq��q����ͤ����oWJ�f�N20~V�Ogr/m��־"��qW=��� ��=����l����PYZ݀C2c�*X�y�GRп�v.�Y�/U_� B61Ho�h�|�0@xv�XmC����k�����q����j./��{]�-g��,��4�n@_#vjΚ���:f����}�C��ϣ�ܳ��)�I^��L��������'!�{��kx`�(,!�=M	� tQ�>
��Ē4*2�����	�g2>�}��O%唭�c@��?�K�C�B
�`℉[�TM���H��i��0�Y	k��ӑk��y��=����[��TXJs`�"�[�܆���:�]2/^����8�v��au�gE�X1h睳T�8E�+�������Nz�W�v<�83)���N%Yn��j����#����\ǵ/�,LrzL�~��R6uh��d�B$u�mF]W��`��j�c��t���P��S�o��Gǖq�������v���4�6c6g�C4ʑH���� �u�	�JB��̻�O��ͮ-�Yj�����RYВ�n�ep_��B�[�Oro��>�9�z���2A�C����{�T��<�^%rY6��>�C�z�K�$fe}�)�fu^I}JȻʈq�(�@*��Ì<����!���M)��4=�G
&p \l\�W3�Aj��� N*�܁�-�қ�j��|���1��m�]@S�S�W?��Np�ݗ�^�sn	�9V�����8���&^�LR�W��;�����o*���Ƣ��+�W�h�������:�N�\���f�C�ܤ���f}�o>����7������Z"~7l�^�K~עE܄Ӥ�N)� �����-}#8�+�6Λo�E7�vV���w�y5�JnF�� ��
Q�\���w3&�@\�,//SR��+r����J��)HA���kN�	���ij�z�0�J�Y_0Sǚ}�2�1���H?SleQ4�Z���O�w��O"�}��.�rwc�A���-p�T�ĩ�k�QT����Om��;���3e֦�뵛�O��$�&��'~Z�����J�,;�>T����!�eڐ�m?��< V��*�$2��E`ա������eNng<ҥ�c�e$ ��Օܝ��r�)b��@�$�q��$DC�{l�l�( �Sk�f�p?�*,$6x�q�4`�m6���jq��x��j�����Q�h��s��]:�=!RƖg;����l�����d���j"
B=���{�>K�<���*�gSxa�n�>�%�iT�����n����K��Q��u�)�^�jg� S��u��	��)gD�9��ϓ<��� K�T���%x�u�r'q�M�P���q#��W�|��I��B6�*��bͱ٤�%�D��oK�JcZ�D^S�
�-V�h��F������5g��C�C���XG!"���3�v��r�11I�$��-z}����ɲy���L7��B�%��4���Z/U�g&fM��x����{�<w�ƽq�X	(����d�tH��q>ӯ��s� 2�ʘD�SBX��π���ł�Pz�~�^�o4�#P��X �f����M=!!�?p_��Lz���6��b��Z�?�͢a�<o(I�Xv^p�W��h#p�&Mr窲�X�0ŐV�	W��O<���>z�D�)���<�W�����	�`� ɸ�na��0�ω���9U�-���u�8���Ä$�������	��o��~�l�d����XER��a7��f����B���r׻�� 0�G��1�,P႞	nW�.=�\��m�Ϣ�.2�&O�%fo�y��9(��9H͙��� ��:Th�9 F��
A�ԬDyt�vt!���HN7��Q!Q���-��Bq�T-#��!�e�
�*>+ekJq.��*H-�������z�X�$h�`�q�Aq�^Y����,8��9i�#�l� �#�W{OH:��;�U�"�!��������s,�v(X|�I
�dށTT���M�9���s<:(��~co�*�GF� �p��#T��4���k<z�G�u��K��FɈ�r�ʭz��m��aDD6�U{\3V�Ƈ?(#�1_���x!�:_������k����|�ѡ����8���7�&WW�t�њ�t=��k���q���9(?rv�\$s���-��9�xqQ#V�Qm�2 ߁Lǅ��1'ű�m�	�u�������=���?V%|��n�aD:6�]~?����$����4^so��j揦m�AyQ����6>��-���O���'���_4���͒s��|mOk�{ܖ<��D��Cb�+��}/,���\�s!�?^6O����bP!���'��1�X���αl�'�Z�`/��*�1w5J>aHsܦ�`]�.Y��N��R<��	��j��)�
mba���"���Ve��:��7f@�,� ��˰"��=��I1���4�x��7U�O�ޭo��R�C���ỹ�՟ܤL��]�Pau��y��lJ�^�G�^F>^2�\�=\������z��%Gdb
ݔr�a����,xR�c߱����ßDzS��)'�?��`,j`�4� o;��/�˂�y	�í��y����[R�o�K=譧��c��x�����-.��TuN_Lԧ��Su[�v��燧+4�_q��Ot�R+�e}�b�� b��V^Zx��1���<.5ٰ�
-�yR ��KL��!���M�W��v[�K�'���@�1)1,�R�^ci����*��Q=�\�	�Y��M�"E��>�ǝ͞1@iw�-|y���X )�7�Cf=�:���iQm�6�Q��\B.�l̜af���c��7����A���rp�7*Y��7/��M�.J�D����%w���RgC4Jt�=>���z��\�m��fL���`C�N�ε}�+w�I,AD.���%�=l���aS�*���1���5C��C�{GmM�h����}�V�'8�hz��J�StۤQ��'mG�L�(7�PYs�L�WA,G��F�Y��ڙG�7�g�&�j�"%Rq�~,�t�Z����t���b�)"�����B�h������uׯ�����L�[���1a��e�{0�)��>pp��ם�g����3B��<���=M
_[94�}�<R�g-@\造�Kٚ+�_��C��d��櫼UU&��)'hU������
њȆ�{����[��s����]W,���f�˝���2o�O>�S�4l�c��M�E�()ɲ��,���7�9�s�����9�WH��%dg[�rFO^�1���s����c�HJEb�i*k��R�eeh{��1�SCzq��M&d���,ֶ�M�$w-\��Ju�k��<��c�)��n����e�3��T�w�}9BA�SBKRcP��������E3���*�^��d��&��׌T�H�R֎i�F�X8�6٦��L*���M���gM��N��P�A�E��u�]Ū�Jz���32,O���m�k �T�
8�bx~�Kp��&�/ �q�AK�P+b�&���s#��;(`�S��pO2�����Ȩ������j��\+�c���j����v$Xt��y�Լ�K���#Q�$4�{��k�r�-�m���\W�4Xl�6R��(1�'����.��&#"Ua� ���{���Mr.0o/�0���3p��'�q'�z�A�P���:���E�a��e�O��g�ih���wUZ2\G8Z
/�\��� �p�7����F4�5�jK${Ђ,;T�)yWܥ�b���%x�m��{P���U����ћq�R�7�-������P�$��1��?B�3�"rF������cD~ۖ�[�@�2$M;��nH�}��>1�֕>�i'�fd���M���S�Hݟ`�?/�F_��V���c�"?���:��hUyeg�2���A�B��5�F��zi��Ԕ@�{Csԣ��Տ�?'�BX_�!����c��DAVh�r�w_Uy�}�q�R�Xk�/�}��YYl軔L��& V0_1��s�"�Z(q�x�Z�y�a�ͪ�/T�Z�B��l��rvW�c{��i�P��l��;�5[�s'��I�7�X����9n14kA��!6�kB� ���Aȭn�҈]��E�30 ���۵LT.v>_u��JeQ��@�ƚ"u6n�Ȓ�y��޳���n���q�5G�_͜��F���Ӕ��:5���<<���;&Y�&׌b������y�L�аφ;�v���ѻS��=�4����9e�[F3���{�ZWVK� ���"S����(�Ez=��e�C��˱#\΄P�-	ahs�,6����p�׬J��.]�/N��Kez�b�܆��~F8#`B�Κ�9� �\s(�mvZS��U�XK^a����@�dj�8��ɺ�\�;3��	b�˵U��S�{]��À��*�]���#	P\0%ʡ0�d����m�{;AJ
�� ���[�m����ٚ��q�I����_�H8~��aȵ+Ŗ�O��~���i��
�HJsl4���s֩gh���p����=�W�˭E�1ڧA1��cy=(��.Z�s�=8i�99��(��jt���⼩�݁� �� r�V�9����oIZ���*8��E�QS�b;������SŌ�� ����&�՟z�\�C91��4�Y��|�w`�]�Mߪ��q�:+fbuJ(��B�A"m�J�֕!�Jmi���,W�zKT!@�ȅ��|�j�86�<3�Z����C�q�����!3,4"͈�?,�ӊ�x��C��?�;]'���j�}/�L��ۈP®�V��?���\L8o�t�.$��x���`&�N�m�F��nCt
`.�{\�@''D���|�9�Q�捽�<�C��H��'�P�}�ZI�ĀWرŵ���:���k%��t���ϭH/�l�H3p�o��6_tf�ɀ#���,��馎�7�3=GG�\��kӉNc�aV�8���΄-)9�ׁ��6X��@f!q��SK4�षB0��2��koC������.K?b��8�~k�����x�U�]��m4����)eͨ��~_￝�}C�J�>�~�/�C��?�WWt�x���Cn,��-7����r���%�L���Ҭ{Ѻ�d6w���)ܾ���8����[�|[��7�~pA�NR,6W�C���ب1�ă�v�ם�>=��M;+䧱����;%��_�g�3b���9CW�m�@�"�d�2����|�o١�g��g��r2�Xv��0nN�_l�����)�Щ*U�ldԆ���4�:�%$�T#b�Ǭ�+vM�5\�q�����Ix�d��([}�=y���j�u��D�O'�I�RDˉ� ������J�W�
2z���_��_�7z�����0���貂�wdN�ֹ׽����ݬ'��O���>�Oa���Į�}�S݉+����b�/�׽���$���IˢS�P��'�7�y���3Ҟ≒]F��ړ^�zmys�c����`�,�נ�
�>eH�g��`�Fj�Db�S�1�03����c}v��
�=_x>�K
�:6F��:���x���u:8����Ѽ�I��W} ���L����i`n���
둟���4�ߏ��讏F�f�}y$��t��5���@� ��*!`�����W-�α�<���)��MD�b��图��G~R�����E�l�����_0.���2E��-5��{%��5�=��q'�&LJ��YaKNI��HLA�������!)� �NJ(`+�N�,MR�,��g���<��X(�T��u(�';����9C��(��5-����i�@���d4�Sl<��9Y�������M���@
"�e�&6��m����Ӆ�1	ړ�݂K+�C�Avѝ���s��{'�T�#��;H��^2��V?kĻ�}pUR�D�N�	�!�V��,Ħ|�&����>��͢Y���X6H$D��$��|q��B�G�ҙlk��N~�t���"�>�H�9o#�����8��Q�n�|'I]#͞�I�q¾��fƱκ_2��M�*M�?�grT�K��a��֘v�$�B#D�@�뼓K-6�B8]�����~:�L/���c �J�1�8!e<�[\m��/??�`M�< Ȓ�R{�&* �ju�k��!]:���e�"բWGZ+�t���r��9���ݪZ@1�ZwE�9eضg\QG���-Y0m ��ѯ�ܳ�n`��C	KWyV���ޛ�]�ˊXZe���`PD��R%�<'��d^p9q8g���u�����܎��Z�<T1�ޚ��$Be�������S�v��wX]�9��?{H�P z�}=`Ir��+e��V`-X!#�ŗYޛ���>`�0%�{�_>���2� >�]�'T?[��}7vxδ���l�3�m�o"�~p�m?����/�����Ʃ]���|	�Y��O�=b-��ih��ӏs�
�,�yd�=Y؝�I"x�]�S�zy��z�]<&�q�Vk"���☗,�K��1"K�c�ˁ1���]5�R���<y�$�-��g�Ԣ�~@�@���<���Ft���'���r܉�Bh���}��;:Z8�ZLx^K�����O�]��QA�W�`c�s�Ϯ�|T��^�<�׀!<�5�Y;b�^XK9�����5�
����(ɓ����N�Z�J���ݢ����{ﴫ;M��������ez�IU�C�1x���ynܚxa�W��1	L}�}��&}��h�JMM�C���u�6�:��0.�~���&���Z0 ��EF.�J��ǰ_�Dđ�M�U��Ma�sK�H.(���B���ת�=������k=񆮪#�߲�D�Xw�]-����w�nVK6)��5��L3�8:h��D1`�� �|{v�n`]u�Wk[�J�:n|��%�
�mR����)aFR$$�H�+�dԀ�o4�8�r��f��={�T:���WR��c�E��d%R�,�m��}K���M�_qcv�8�T�3Z���&�+�(�P��N�D5�}��cyp����z!����o��ILFt�Ď�xV���L�����6��96! ��r#x) �ŋ�o��J�UL-��wV���Hg��U��_l��^<���E �k����Tf)i{u�p�A�ކ�����*���lAT�d���F��@ű�^>�IM���pC{$�����=+~i��X-Q�Hc/>vUf>Ix��M����9�[��V���栰2�ʠ�T�UPN]-7��p���r���b9�c��7�P���~Q2���t���>����C'~4Go �HS���IU��&������B �VZ듃Z�G�hjf��_���I}�Ӡ�D��V?���w��U���^i/Wn1��+6�	�Î��_�� `���?koZ���k�W9�G�:�i�뇫T�	��STr��ݏ�����zbX�C�(tt����Z��EE-ĳ}r{�׫��Wj�.]��(3�PV(`	wh�~�s����(�>���C��[����SlU@���$��4�?�m�q�5*�`��2���|����f�l�j9ks��I�mz�nn�W���W��v����d�ZX5p�O0|�}v�����(���qI��t�@��2:��Y�J���Y�) 8qq ��s��e[ ���Y��:�?��fϥ���֐ƃЂ��/�OCi�6�3ХQ���U��£��L�.����UcqG��ze��C��"�� ���.�%�!��(��>=����4sI�|�Œ��^�P���#�h�n��6ڹ��V��C��S�q簸4��?�ydM��T�
�r��S�Y��r�#h:�;as�3�x[;i�(|���)G��g�!+�Ѹ�ϔ���qHK)X������� $ўY�އ��UU}�@Y�a,�o�X4(�d`ԡ����mGgE�����a�h\�B��+G?�s �D�� ��@�� �g��M��3��ҧR�j9�k'g,�"��r�A⤚`�ӫ��>q��@r���P�:'�U#��_ �AZ� m��@�@w����o�V�Ɋ�:'߇�<$�U��w�F��?[��Q��Ȩ��&�}�Q�d�+��� 
w'`Cs_�j�Cw���m�X��K&��R9j�j�yK�mz���9�=R�m���F:��	l��9fAz�2��_FF&����Z<RZK#	V��+HA)��cV�������1��s�c������{4�I�S�ǭ=��K�3h��^koKy��_H2�(�׸��X�見�p����Ň��<�&�5�T����E�[\��\~赯�NuhD���L�k�{�"CuS��wOQ�������.c���)ا�i��D{ZZ�{&�=���rB����mo����٪�f'����g�q�*}K1�2��.�Xa�����L3T$d]>��ۂ�Y����9Dlm1.D��஝u;�~�3�Hrԍ67�=����h�=mQ�i�N�����֩��[��ü�p��vi�m���FQ�9���DC[8R��$��2S�����a'��P���&q�x8p�r�r��W9�x��K6hN�+4����0:���ы�?r�1��k�D��܈���ln 	D�v#��Z��V� ���Tb�a���9{@ߑ � ���"a9nG�� q~�Za�R�d2�:7�R6� "f��w��\v��eW�E��ߠL�z�Q�6�x��T0#��D���N�5hꛧk�k��z]�	�@��KZ�T�>꾘���khx�u�>k��e �ޞ{R)zz�}0��-aZ����4\�Ak�[���g���0���8�Xf��B��e=Y�j �e��TxA&O续�a�O�D�O�YDv�%��D~�+놰���
���=��׋z�Z-�6�޲�T�{Yp�]+LF@����׌���{>{��v6�	!�+%����5�F����h�(:��g_��ڹt�!�UkP��r9v����]�m����Hp9n��cهV��� �A�	Y袎�r�J7��M�=!"�L��7[;:/�H���m�n��a?����	B�ܞ��M1�Jdڃ1.���6���u_�;���ZRqֳ"��3�B�Ih�����%�~�!�%�nl�8��<oz��T��y�Ա�I���=�4�}���df���U��*;����)�k���;��關a�ߖ-���`�V0Z��yi��R���d鍆�� If[��%]���y`B�d��2;j��(�z�B�Rx5Waa�C��E���d�:쓽��槕Mw?g@x&\��l����X�9��Y�n�f�Ձh(���`�_$�#��r1ؼ+��I��1L������8ݼ���oWt���AV��LM�3VT6{�.�*��K�K�cU�f�3����w�L)�/0�-��h�����"��@� ��12��[YM�7Zyi
آ(����y�n�h9C��">`�뙃�����é�u���$Q8�dQX��4Mg���b��1��[Ø�sZ��7��^��,x�7&6�����17je��E�r�nX|!7���{�����ĥ��������6b�W��[s,�v�`���+5��/���.za�$w�,�s����/���Г0횒z�J)A��8V�Q��u)g9������A�+Hm�����ߚ��YJ��!��y���f&�iP���r��%5�,�")(@ŏ����^��ᣦ�)��4��nU�
{
F�D"���<ڊ�ژ�]���4}�Pp��c�n&�����:m�gj���t�4�8�OJǈu�l������ �|�Mθ̢0�O�)�z��E����M�Ɏ�*w�����o��p�hNȺ5��N�H^=C����]�S�j8&�{�Ԙ�J��?�����Wb�
����<�T��t�.��^b�T���{�y7W�u4[��{Ô�;0
�;4:��=��^�x�ܟ�B�֮n���1��'�xt�85M�n�`�e���GU't.�1��/�/��i�(�榚ڵ��-��w��n�H������'蚉}]]�F���
�.�1|f=<�
#�)(,�/�?[Xib��-7b�����&jm�����6}@}Vf#����^,��+� �^"x��Gޔo��)6����׋,���E'5� 8z�9�7Ç��<�P3�f����Z�i45�%�\�j�E�(��D�
���
�k���y��nRYL�u4RIDt��eS�,8�4��,�Z�RSd׷6�Ͼ�W���	Q9�9˛\��>V�{�錗sw����E�k�0��2���=!��t�#�U'�����������ecb��x��G6@������f:�~��4�M��#wo)�>��S��$a�z�i��f"��"w��I�U��I+䡎��*��i�޼c��a%�l�T�^W#�@cU��~�V̚�t7��F���z)zU�{id�H�+>�Ҝ�	i����?[m��WF���9d
�5����}�Rx\(��B_�\e8�ix�R4I�Cu���b,Wu��/��������ܰ?H.M�G�u�L;����ۻ4�.�FC�˻�>��#��)�!�v#�K/}���;q�}�z��Sb0��Z�����(�����de����Z�&�)�>�P�98�`
�0��;HR�J;ȢєS��m�2�
N�/�b��7w�k��)>���e��yF�3��J�X�H8o)�Ml���i���~X㍑P	� �:P��TT"V#2nl�_��Xˆ��D��V&)6�4~��)q��h/=a���y�=�bH�ŸbL�''a�j`�o&�2|�,�ksl�u�Hӗ�axîK`����}.,�.~��ٿ�C7(6�w[�5v,E&�߉S^�CE��ى�����'?�������A�eY�Ǫw�͔!M��>Ɂ�:�?45aދx@��kAU��P�B�V�p��6�9�X���Ԩ��R����B�P�4�TlRA�AK�Q�RxZ#�k�d�N���`�I�rˊBz���}JY��)B]��!�s~	�xbo$;4������:h�0*�j$FK&����}OÀ/Օ2
�Sp��hM~\"w�I,f��m�"aYJ��ES� �w�e�'�6��q���ܱ�H������ݳ�-Ј_��)�<feO=	��wqxjk_�L,y��A#S�>�l&hT���OVة��>9�Wݻ �$�t��G�`��H��E-�a,*���K�x��[M�ǈ�].�Nu�T����Ɗ�Yb�y�:^@�kJl-N"��=V �zͪK.R�9�}6����ͩ�/K�
h��a �f?�N�ǎ�{�Ҍq%�cų���s�OvL��tEsx�5!|���p�|{Kf��ɏ��w5�=h��#"�$�뫎���:�fR�k�P��D�&_��NDL�)��O����=����r}��)�u��D�r�Iy9�헬4����F~8 ���V��K3��N��UR4G��2�6�Gd3�¦�PZ剃R{x�@�x�p���U?��yq�}u-֝ B��^��U�%��
ڝZ�
V^j��@@(kJ��v-��عU��2{?"�VU=��́A����)��)[xS��ٽ[��x_��.�#�zq�);\��w6��l�Ua���w"����&+D�m������Bi���OĨ�w�K���E6 y��i��y��uփ��Ň5J���^�S��	���}��Q���+����}���|�TnKQB�z��|^*�*��b#�B����܀�7�re��9H��63��b4��R���I�n�"�U�/3:�Fа`kOb`	冡�?��w�6��/�4��G#�6�߬� �P!2<@���Cp�1�D��߮������;�IWgv�;�����؋\0�lO�p�0.͐�z��t�j��RG����)���?�9ݶx.וu8,�2[������ă�lԧ�)&P�U0}�s�pވ�8������h�Z�JP��^��D�p�Ya�[�Ӊ6S���kz~݊bڈa�,���vj�j�u�_K ��h8<���j\@^�7@h����������4{�`ȵ"� bB���B�'0�J�	�T�;�ˮ[����Q�(/%n�d�O�x5�za
X�}141I�E�z#_F�sl���>?�'0/��v�V�/���đD��x�#��c�������v6���nN��{L'v��KM�I������E)���ރթJ~H����o�����b��H��
=��P;��g_�D5���{ٔ���㽎�z���W�ɻ
t�E<W=�Č=%q�{������&�b+)A�Fo�=�uݚ�k]�	�d<�Yz�O(Q�ʭ�����V!6EcO�� �FPDi�&�~�G��sOk,�#.J���,VcT����:�u�Qsb~���ܶr�~�\C��L�M4���yM�]�[d�ϟa-E^Fŵs�Y��+V���R޷�"mZ�)�Ւ�ƍ�i��0 �-�����ϻy�
fXy,�f}�p���#����e�Cޫ���J4�1�9�T|Ɂ�*���J�0����������������m!E!W'|��Ǖ��9h��p�13�z�د�t|DHB�~���t�����@F`���F�zW��`�83���:�7\VK��̨Ԯ�+@-���Z�f�?t�:���jދ�ܛ2f9�\o~�n�9b�:�$Np5��׋�ȴ�W��Bp� �6�`���bqD>�<
�_�KmǔX1\ŵj:�����Ƣk	~�_z���t~�k�p����'l�:����|�`��q�c��Vț�(b���7b��ӓ��P���z�-n6����Dn�x�#ik��s (��
(n�#�׮,�Im�t�b΁fQ�E��~���8�u��V��r$
xI��M\�8����J�>ƛg�hWZ�Vt�+�O���X��wG�v��l�jҝ�{�����l�|�Q'�Q���Y"�����~S0�Q^O���r6��xD��C�"���5Z�6o*Vog޿����O��G������D�c17i:�b7z�qkL����>�«� �c��p����������I�̀�>�C�����g鷑Eg%N {���(��^�O#a:�TD9����P�R���25�5��M�YJ��^4)���d����G�ѧ��@���&{���d�S��bm����x%���f(c�19�D��|ଔ��PT�vuOD��k9����\�0�?�uou�LR��)���Epv���?0�T���}@"�5��"�>�+�ݸ��u9��Y`*`Ҷ}����f$ׁǏra�ް�Q-��9?z���iƍ?g��Q�R�9}>kT�Hŏg8��m�on-:�����J3V$�d�	�q!<���$��6�i-e<�fh�_1H�Q���65�ը��e~MƓ�.�u�����R�|��:Pk�s�����K���B����<ן2����`!{��)N��`�;��چ`YaϷ٢�����P��vZ�U�#����|���Ϻ�FϐWDf���a�&��g!Yh���u��b�����~2�N$��W�,qr��d���x77�����\_��iB>pq&�Nu7nz���?�Qp�:*�Z!���jI��oϺrZ���:Lwve۬�މ�%����g��`�_�qp�� y�A?��x��V��V?Z�^����]I��c��HLw���g��eK#�˟��������V�ȼ�����2ԧ����X䬴<�(��eV�rMq����'t?�ge�e29ˮ>^"��p�/��o�)����a�����$b݋��;��I�a=�9��q����E��S8<�L|��O댪��j\V�W��I����A�ݖAat�����~A�c"a��.�I� ?���q��&>`���_c㋆ �X���!�N��_l��VټL��}��e���Id��K;;r�i�>iz�%@ƑtJ@Y��B�Be>�>74a�٨�ȯ�{3m��(�0#d�G����&��&=/�B3^�,W)�/$g��p�lw�BA�j����؂�8c��Ce���T�^�K������
˧�2D�� MK+b�0J+tn;�.���Q��CP:eux�S)�Bz-�rL����@� �C����kh}���@ڡ#�r+_���v{[���<d�N�[��p-��XE��K1�0I��^��Φ˗�$O��_�a`�8�Rڡ�^��/�D?e�w��O���Rm�l%0�Yi��E���v�r-�8[ʃ�I<O���0�w�gu���Q��$�@�\ nl���S�X�I���M��;t�X�Н5��s�H=�`����l�B,qPe���w�V^����mq��!U�y�����I>��ɖ�X�b��N)]ލ��W����C��(i�cT	���ۤ�E���aB��[�9��~��U����d��/��%��g=Z��)�dWQ�h!iY
=�U��?�[�,2^�n��}�K�Ccr.K����|�\���H�X��p�w���5��1L��e��H�Znyl��j6_�T�[����n�@�َ~Ҙ<]â�"��ӧ���.B�f*��Q]ֹ��B�ً���֞�p �0�we6�_7�0����� /��j�@2�ׅO�<wN�̷�1�z�ܜ�u(���x2�!V~�'�QBT䶬���/%=�ѵ�T]ը¹%�R�"#-��\�B6��ɓ��u�FX�g$��4;����q��]��%܎|O���ߘC��+�nA��T�@�;�Br�PL�zp=ۄ�	�N���|�MH̍�K�Ȫ,������W�%s�ř
��O���e�靮p�?g�����
S�w��hIEGw�7��3[Tm�Di�9��|y>9�-�Y.kC���-���3䙦�w��:�u�r��F*� L�,��U�CmWv�� th� b+�p��-~�	�x2M&m�FMA�����g�f$,�a�jY^��a�NR����]n��abU͚",9� �:�'X�%!U���f����0�7�!��`���0'�W0
�ﾗr��.�dXRl���<M���D���ٞo���4���OF���Vc�J�'���E ��a��0��O�P-��e��,e��#�OsBN1��P4����6��Z�n݁_5�h�X��A�S���:~ �9Gβ�J!?�\�<���$?C����nl���P-��ϝZ�.xF�
�^w��@D����b���� "�7�}p1j�"�@z��(D����Y��h��(���M{-�N �����\�6�7�7�G� �����U�
��;���s�<_��ս�$|�-C;�aS���S���]d�˽��z����LM�f������%�1]��]0;�X�j���=$��1��pe�so�7��.i�V����h-����*����܋G�-�:[~ͧ �ZV
k���3/Uha.�-Xr�̱װT��v��7��R�ğ��f��d
n��G)ͼ,\2$N��Z$Ȣ��b�;�f�����l0˪�E�u�2�f��7%8�m��v��SZ[��}pw+����d��w:����I�%�v��G;��z�O%v7�m�ؠ3_������S��"�eB��hS��'��'���0��K���#��Z����P�<�`�9x�t���ǜ���nND�:�ǫ������L=���=Ϥ^�"��}i��Pm��(�u�EĤ�\�$�ҕ���?�d`���\�b�Xcl����͙惙ZZ�H��*�-U��-C6�q�7Y�_g�I��In_I��Ԇ~�o V�u�Wn�GB�W<D�?���GT�>���
��'K���e�����*��Z>6�NG�����[)����n�#��&粦�[��{�]�q�����E����X� ��:-�u�z����ۼ���J0琤h�M���.p�/����
�ok5�a$q���v�D��7�"V�4�9��J��g >�u2�b���K:PЮ��Pw��>T �*�Q|�Τ������;fn;���]�b�c��;�|'��4��)�w�q�� �{��[��m�3W!b�]�:�<�U�p��lW�gd�eΆ�6���\��>� y)Xj�ՋM1<�6r��?/�#e~wL�[�
�C(�N���iѨ�2��n���+����w3~r����!3�,�:jSa����I�t�|R�� �%�Ń��!<�K��B���0�xF�q���8D���Z��'ѿ�ʰ����U�c�7�V���(|���T���}�II���bk�[b��xoqUvk�VW�(��[�e�c>�I'��5�o�<
�����Ѯ�B�Hʫ8PO%f���	Ǎ��SH���N��Z�m۹䔱r� TJy���;�����W
n���J7"�ιvЬO�6�Q^�x&�ϭM|gW�y:$�{�D�B�k�r�po�(!�9��3(�n'�L��������,�!?�#49b�쥺��p%Y�&�S�)���>�a���yP ��|���ɥ5&�J�"
�ig��ʭ�m�d4�+�G Q*mcq���W�����p0�:�$���+�rmThS�s��|At��f�$_���: ¼�`tjBxʶ� [ 4`��'���X*��	�E[�Qds�냟;�;xk��9YmGK�{���8��"}J�4�S��~z��t�b����nv���o��F�x�""I��9s�o�H�'���ZS�۳��mbAR9�+�ʭ{h��
ֵ�Z�:�a�ӫ>F��C 8���_Y@�áHg'�ʿ���A�e���;��8B1�� �. ����C��Jg����c�'d�8���yf�ݹ����#4@+�,��i�_q6?�V�u/K.~j6) ��p\���쿇.!7�ud�k��I����,��
�-��jC��%�n���x� $L�6������h�8���|��{ͅݗb/Y�m2Y�C��H���b���i�M�=��Z�.�t�(�)�p������Rtv� �k��v�'7s`B=��?�����?���y���%���g9Ƭ������GF�<�(��J�&e1�*����K%�\ ���PIמ*������.[}�'%��{��9�����n����I<�g/�1�f%�k;ʮ:��~�b�g=iY��x��<�Pʾn|sU]�V��5�NhO�S����� �AU��23Q�n��P�ыQN>m֜��`���F:A���v���t�JJ�.�|} *�6k*%��~ud�k-��Eṿ�'�t��
�~p���-�_waVrOf�<�/��[�EV�a-,�����,[��yH&At��5�t3	�\���(p�g�3�ʡ7�{���b�m�E�V�i;�>�<�|p�4� 籴pu.��i�u�!�8�i�,U�"�'����V3��a��׀��1��T�+,�'���'8��S4|�s�	t=��|����ox$V#U(.�K��?0� 7�_F�0��G�,ޔ���*���W��Q�с����%�5���#����Z �g��^�abĚ�o:?�ub������j��Nێ~��N�Č$����a������0"*+&4}�}m�F4��r��[}F"���Zb��Ow*���Րe������	/��M���XӁ�#0�oy-ç�J͍q��˴F�6�w(*��D����:���;^�1��[	�;s;~�4!UՉ���Z����¨>Ss06�D:w�PL<�p�\���� ��Yxc�~V,�'��lYV~����$��)(�4���ᗫks�J����:vvrnx�MOe�;J��Q(��h��`k�F	�������<�jT@��K �e�A}n%r�S�8�"�@=�#_�I��PȦ�?N�0�C��?��E;`��S����9���
HT��'<�HE�pog(�$V�>��0��������l�DE��j��N����dx������EnT7�x��L@�_��LG�b��=E�Z��3��~�3}����x�?�_�ĥ�6 �.���c��O�X(�$�L�(�<P%b�K/��NNn�É<���ȯ��r��U��6���>Y������v��������3oh�mˆ��+��ִ���g�N�Lo�+�#NS��HT�Y�)�"꫻�3yG%C�$
��lX=+C���j4��R�}�'y�JW��2ƃ�s�e	Q��"�o�x�����8`32�O�?0L�����R�,v��w�u'0Y �
`'���Ώ��!��E�2ا��T��d��ϭ�y)���ix���� o��2d��_����)����
�P�,�}�>S�Y���QP�3Z�N,�5X�5!����D�<��ݩO\w���'$v��Q�#j5��e���N� 0v��ŷ���E��1l\�ɓ���M�S��`��g���r3���
�2�[/��~����*�M��I�b�P�^T	O�5(~}@2�GK��Ka��N�W���K��[��xW��w\�g����$�e��bF7>1;0��Y��ao(l7D����+�v���k&��E.5��P¢W�-���J�X�L)��l�R�0� '1=�����b<����m�H#&�tE�w�=�T�@�Jn�赑����1=2��|��LG��@5�魪G���5b^=�`��H���p�/O��s��R��x��6�KQ�f�I��亃�:��T��9�oܐi���	7W��x;{%_l��ɪ'f��Q:�;>-�>S�&;�$_��B��NE`L�u]ҎN	7�H�[�S��.�MURM��e0�����S�]KW�F�A���K�+N�������۽�N�OPa] �%%=ID�ւ��[u3i�����8f�����B����e�[<w
�_�������q^W���)#R,��P�ݹ��mk`91�vX��y�3��t�����_�s,��0D�J7I���`<Na��|�W&5���P�j�H�Λ������o/wLK���qz�VZ"�����N]��8�����[5����-��Ǟ��\��{M���9NsZ��X�	mF�~��]L"��Z痣!�b2c�n�p,�/�:sQQ���y�q��������\��_W�l��Y؜���i7� ����ju�
�����%J٦��iE�)C���#x��9@C�R����N�޻���qȥ��0�7!:��zNŷu���	-s������왇�7vÓ&h�c`�.**���h+8塘I[�9�`sGS���Mk#������T)�p.��!��;29�2&�C�x��7� ���:h����V����͘�P�u7Vt�,Z��f폦��obZQB��]�*`z2b��2{�)ǡ���_B���ų4�C��3|x 8Lf�,%�Z I_������G%��swM�~��!�$SR؂�c�.���D/Q$�ƀ��H�n��T%U�����dk'��q��%bmH��$�Ur^t�<�"���>���!�;�' P�[�6%�,��4/�(��ϻIB.{�Wd1OS�-�E�\��\P��o��C���Y�HY�cꅼi
��j��o�º8�����8����(>lri|�נJ�/B�P�Lb�s��a���J�X��9Ȟ��)�6)JR��ڄ���k���8��P}��``)�a*���Kw>Px,��)��s읡C�Z�t�����=	JI�b��|_ QS�CF�H'hj�0'�]׀w�>c��B����~�о��g=�G9�W����M�s��\z�Hq�f�46��͕�X�7�<�oc�)�ߠn��Ԟ�u�qV�Ƴmv�"��> �Z�!��aMM-No|�c��	"hӁK�N��*{�hSF.�$ԗ��Gg4��	�n+�>Vv�=�f]���m:h�FK>����.ե[�$,g��i��-1tH9�8�j!���9���K�a����5M���L�^�4&1����K�>yĆG��i�yћ��d�×�Z�ʣ�[W{L�Cvi�\S_n�@��H�s��z�������TYr[�{z�u�C�]�Gh��1�������F��T�݆wwM�-ֿxu?!\��.ݪQԌ�~l����%?hg ����,'<L^/�ŝ�5U�K�"�d����/mzr�&#+��W+�+�1�6]��b��<�q�us�Ԫhe}t�[E����0h^\�u ��ۙ����nv��SK�䭜��E�^I%��l�.E��=�+�i�w��}��%��P��,��h��@m8?iR� �����\>M}�4R���L��v���JϤ�����G�s�s�+(6L�%�Om�B�.�sP#-�%(����4j���V~�������L��'zc�ײ-�-�/�k7��N�]z�| < V��/��zP�Q8ky�ꑷJe� b�.��s8$^��Z��Љ��/�,�+!�D�7R%Y��V��
y�ѯ�����G�m�9�<��>HgN�}�❝D3�̕G����d�a��͕ny;z>�%Q�G�;���B�!��c6��,�!ђ
����FV4��*��."�>1 ��4�rAӮ�n��!�g�[�с�a������"��h��A�BQMy7YIN
tX�5jy�}��2t��%�aF	�,��2m�>q �4eyܧ-~��� \ ��I�$�� i<r��y����1��8)�3����Nl��0�>�#��x�6���*�2���2������6+�<�:D\�J�S�VTq-X������<nZC���������
�μ� Q -��_���jr��2T�Ƽ�w*�����/���@c2O)��*&���}�[t�ڤ�7Wq���r;�ߙc�:�_0�C�W���>��l��?�jdd�24H��'�Pj	f��bIX�Wʔpfs��0�9���>�7�#����a�DոZ/�*Fs�� $'R��\Aۉ��J���3Z��МE\/w�~���z���[�߇֏�+ޙ����h�I��4]R��;FM��8mm�̝�$����F'8�NxG��s#ݎk?%���Y~KH,����q(z��#,�n�++� �:�b������p�����G�w^�&��9P��G�C��\Ә�n��'!�"6�,�z��{
�lEF��X���<��H�����F~O��[�ڗ���kX� 2���ÞT�9q��������D������b�
�u��C��]��,i+爩N�ή��6�|φ&�E�"���Ȉ�ч��utA�:��L� �I����~2i})��2��o�;�L��
b�b���O�J�۶c�~��c��j@<���#��ʙ"�԰s�c�^���V�P��"��E
�?x���ݲYb����)�$O�ya�t&��6"�'. �j� -\�/�(�0W�S�Tn2��G��q/��5T� Fc|﵅���5�hA)�� )h�l5,&Wl��i�8R����W�6���2��0�0wn��F0����.��[S����G챖�8#�[���H4��IfHqz��½m�zl�)|:h�l1�k�7$�6[{��͞�«*��Z
�y������.z�(#��C7� �G���T&ul��U������i!�Db�*a<�����/t�Ja��c.2D�9��?}��ɺ��ܺ� Ҵ��	%��eSv��֬������盎95E=<�x]�?���}���#g�`�|��^@��O�$�YO����yۈ8;މ�]�0����5%��lcl�Y�}����ŉ0�ߚj�R��]y!�׎G����dE�X-�6����{ُ"��Yz
o~�����Q�z$�i�WT���b���#(2�Y,�߭�e���-��L��m�`b��JI�%���90�Zd):�����rT':�x�I���9� !�!�e�ޘ����^X��C1Ī�9+�����Ȍ���/9�)\*����(_�N��.��������T�n�M�V"3�/.vGG�p۴��^ey�a=U�hq���^ݴu����_��{X����)�ʣ�8*�TNN���d�����4��C0-�G�wvT������#����d��z���6��m	һ�~C���ÐA񠪏_*������l*r򛺒��wo`�Ʉѧ�����jn�0�Ls ˇ�vZwm�6�ۆ�:�F�RŚ��{*�,97^���4{���j�ȭL�z��@ɸWWz켚�4�����9��>�����i�䣪�L�o3_A��M��0C���	<{���+����\�L�u�/��5�#P)��w���n!�l�Q,�x�'6A� ܓHL���ʼ����r��|���)��U˕̗����L�ҕ��pX��u\�Z�/o?�|)�D�O
|ߢv}�����썄��}��}�-HsLOY�}c�j�J�a�����s7�����J~��:�F�=�3�x�QX�W�c����3=t��Z�Ӟ���n�{�9�4�/�/����a�(�w�!`<z���;#�J�ӗR���q��O�m�q�i��� ��]��q[��*�ӌa���RK�k>uRmp(�=���۰������qa5�w�3y';�tt`��E_�i��ЙV�3֑��Q6튱OT̜/˪�����f�:t"PLgw���$W�l=rq:���Sz�yщ2R{�~����i	$��mB��ܐ�A�id�G��ὺ��t�ezf'lA�����30@����ֶ��@�o��2@�XP�AOO.��Ċ�-~�q�ų��$�F$Y�UYn�(��?YQU�I�p_>�϶�f��4��$̸��q�P_7�>;�*ec���.� ��Z��^��I�u�WB)�#?��
�aV�[�$�i	�D�M�.��ЉW��.c�Y��B���LC<5�$dC?��$ɧl�� f������
�9���S�o溽�c��T� ��@���W���P��+��0�zda�IɝP����0��ݢ�tHR��z����	�^4<��^��{{h�T���Y]=����c�u�"x���x���G�g�7ѫ��U��4:)�Q��؇���>~�c���,��Ǚ����_¬��yCxJ ��M�5%��2�����=JR����B�7d��%O���ç�r���I�4�\G��Y�4�E��	7�gk��<���	`Gۓ1�+�)�}���䧳���B�-4;�X�]:dR��q�)n��:C�,u�� QB�UQ~ÍZ��D>�OCut/��-nl]$1W{9�hI.�x�X5�6�a���ⳜF\n}Lf:���\=�����`jnAy�PT��bp�� ƨ�7Z��h ��!Y!9]����I���:�eӿ�v��Z|��^�}1X��}b�))K��`��@L���T��}-0����I�2� 	9���<F�J�c2�P}�~�_Tt;�ڬ�u``]�,�Rub"��!i�ٝ��Lܜb7,�|�Ϛ1;g�)��݋V��|}���|�Q]	*���Okml��1�J��'H  �P��8��;�[\'[=xzt�����T��露w�#hn��j�g��񶈩���ɼc`o*�ፔp���G����1�̚ �cA9�J�2l�����L�Wr�&�s�ED��>�����6�Ɍ��D��f�t\ӕn�d��:_�wX�Ќ�b��X�v|(���#[�P>�(����,G�7}��G���,���l��yP"=$;A���a��TG���.'�uH���A��Jk&é�ɰ�:�%cݶ���?L����$�+����ж��S�Z�M�5�|���\%�&�P D�OPZ;�^vWx���>����0D� z-���\U�����4uv��^��
�sn�O|�Ls9���p�����辷̧h6P�}��2��y,c.����?m�
����@-���Pb�QD��P�s\�m(�~y��+�%��ٽ#�ȲSN=�=�Y��1'� 4ٟ����b3��Hڱ"�_(��s�Xyu.�Z�Q��q./W�}H��ke���!#���vɯ���C�����ͤ"��'IK^vYؑ�dl�^�UXE���F}Kұ�oFw�%`yj�Mo p�p��~j�����˧6=�����P����@�x��@n�8��qFC^wy�.-Z.9NO��1���	�8E�сu�$bx*��Q�f�c��3v����
�+�5�D0G���Y��'��
��Э5���î�o�����\͑i�__W�]@y,#НI(��[o���et<�qh�"E�6o?��}�G���V�I�Y[3-��W�M0r�-ڐX��<��Ǹ<c�������Sqw�����p��8�7k���3�bb��*��2̸�#J�wұ.��FMJ���E��9>�?~��j���ZIP~W~��ƿs�i��q��p�V�邎�n��a����8$mE%t$
�E�\���x����c"�^X���b?v�VqX�0?����t����?��Y%���y�A>P��N�]���;�i2�w�WL;4n�
������;A�C�Q*�	����Om�.DH-Ko��Sˊc;!��Lc�!6zF��/�.	���U�_aC��W ��+g�_�:Q�=�7�וx�"ku�.�SR�1I��Z8��!��ў2��֝������S?p����m|R���SgW+m÷�5�f\3f���Gb�����]d�M�ms{��_��Ҟ��G��ݡ�nX
�z9.9�c����dy��.pq~�Tټ�ͫ���+Eq�0�&_e���ɷ�%�ÎW�i�(�d��a*6�FE�%sd����[q����4b�:�8��ơ�\�l������ٗ��Yŝ�l��v�M�̮�*[R%�kd�Q�U� ����7q� F��<H�<-j��|=P��9ӽ�UW0���G��W@���0�A�=�B�ݖy�~��Y٬�W ����"�������9V�����|�W��C-���ԡ����mQ�����E�_UN
��UO?�Έ`_3���-]�љ�B�crCBMv�zL.�Dxk���)�������cw?H��@6����i1�0��E1��6��\��#��3c������J4��� ��B��T�18�$���Kݫ/e~�p��T"�����N�Q@\,֑���p���jb�PB�m�/�u8|_�ݢ.�*��}��;�(����m�ӹtp9G`l,Y��3O�0y�'�j���	M#L�Z>�B��Ͻ'�;��|�#l�3���y�4=�~20�c�FW��3v��J���1�r>��T���T	��U$b�������8ڇ��
��y�U���x1���Ӝ�Pi����,U��!Hih�.�~�����7�"���Y~�����JnE��Wn1�
,^�e������Kf뢙�Ѯ���l-߿�-~?MK�^�m�ߪ�XH�=�.̒��S$M�X쇘��n�4J��!*���Qx�_h���%�{�5)���)���1�TP���n�-�-�{`�_���(�G�TP++�dm!�e������d�F�p;(>7�[�,���)<����N��Yz�'Q\ݚ�yP�t{H��r��&�_N�)�V��.�(��5T��c�)�e��0C�e���)L-�.�u=�"%�}�>�҇�PZ�/�\ir��a��!����	0����/�bF�`7�Uw�!?�,>�d�$��;�S졃P4��+��R$�����§��7��u�Դ|���4�Y�g� �9�����x�3�.Q���G3�ǯ�7�93-�J3ޚR
@'�j �J�U��Ze�@E�P����:�N�f�W_��&4�b����!�K�N� 
?tP�	�&�������9襧�?���T2%�a-�A
8�d{EP�AuN�l���ұ�ѥ�3"�=٦���9�rq!��;T��$�F���o�.�F�{fYV�Bǯ�ܔw�"89�^4�9)�
�f��)�3 �wM�3��֭��G�!��(��>'���|��Y�S��PM��v�DC����(�1.�7���p;�5��;�a�� @խ!4hG�* 2��g�@��ƛ>� ���/���t`��X�������l���a�! �H3��
j�C�x�O\�VJpI�̀X�Od��}A)�:DRBBʧ���ϛ?3��N]=%R��`�5fr�c�?&.�;����ؖ���w3$(�7�c��I�����3����S�n[���v�|���PfU���qI�q��q��m0fH�NA�}M�i���`g���$�f����c3Nb�۞!poXQ���MH���sŲ�Jc4�0+@�8Ƙ���ie��������^�U���7��ط�����-������f^���*�|��N�W2<����Ͱ-��\�J�Ma�os���!�2_)���K��Z�/�?i��2���i�[�T=��E��q
bG��l�J�y:�=o������3�z�"��Ne�ޣ���#9:�-_�<yL��!��N��-���G�0�M�#��6$�N��&8�H���yh��g�jDGf���L��;�f�D��d��	z��F|��y�}&I*W!�!������Rd���[��Y�� �> �H/&qOo���$jM3B��)�&�`�s� �O}�cG/N淙��_��@������s�s��r�q�:Hx���\��>n�������Z���h��el��������W�����#�WD�OEu��
ɯ�2:�vT���G��0�(;�{W�t`/��#���y)�~Oٽv�j
I���}����`6�&+��M5^��a(=�.77�Y��b��CF�l�^B��t��P􍽛S��	��+?t�e1/�.F'�k>֒A�_�110�^+E/��%}k{�<�^��+�;�������WjPF���, N�MkЮ��OE���B K��;�L���������O��$�iZ�Hu�E�¢��KM�f7�&݀
��[�f�]�M^+{�
�%Qm��G��N�DO�|����-�Y��b�������@v��r^�w�}-�<�w��9��8ӹ�Pj#����	Ƒ�_	�*Ę�3�)>�[Pi�P�4:M;u��X��PI��E��r�栫�z0�W�g����٢�߼�=_��oP�x;·8�+��R��S,��m����>A��	���غfǥ�MG�>�>N|����S3XH������:� ��KL��{��Aa�z�ad��<t/(��=*��>ALMZ��Q=��������;)L��5�ǽ��NT��D	��q�&�v��&n��%���j�!l߂E��P�T=n��z%���uҌ9�uEK%	y`ː_�=՜y8� qp���u�Zk��Ǟ����i�Tt40~�F��J����w��{D�kH��;"V11���C\
Y���U.���6W&|&���������'^��|�s�^��l�Z�iT��H�s�E�`y�`��w�`�D��q�٪Vn�ⰴ�YEΕ#�Qd����b/�1��kM+�ʐ~`�����j����+\�s��@�ob��j��iS��Z?�s�Ŵ⟕cf���a� �F��g�g�Fj;��5�Գr`Z�������E\P*ʕ�,%��^�X��ws�x��>|F��A�^���z�Y�D?`�9�Z�����%�mk$������V/M��f]�-�]9N�?��l�>�j�Ln�8�1���ak�� &L
����4�����+x���.s�HǺ@����{!Ί����s�=�^�ֈ���A3��7�nG�u@$
���SE
�K�3�QW����l�0O���	L�	�_�H�/���/�Y�rE���lč�8�2G7����(�	,�ur3�"c6.<���D�����HBAn��zTB>�p�r��ם�v���婈�v ��ԉN��>����
��s��L��)�(|�����(�,Yo3���0#��m �	�U�OB*�^���e���R�g��K'yt�X�@n�����wk[��ΙL� d�j��-�=�����:Gz����
��~B��:4B�T�()���1�M�*-���G�|���Jpx;`(�#[�,sԢOِR0�]�4�؁FVП��-�ǆX-���h�j0[��
l䊰 �Х-Q�գ�̅�r��� q�*t�B;2����Tn�,16I��"I8<I��ȟ�v�[%�Jt��V�1�׉����m1��������Q�!��x>�P#��_�>�<"s�p��ŋ��&37��r�{� y'����r�֠�+ԞhVX���
���G���}��u��A+�%C��M�6�O��Xn =@Y'ߛ�`������Зr�I���gD���=��ɾe��R�"�d�#�59�R	^`)-�E��y��+&��Q�k�������l��|�7O/ ���r
az`3��T��"�؄��| ʾ�n������̄�E(��J Z������ݨ+�}�kC˩�:�����|��a/��*X�]E�x`��!9]^��ۏ �؟�*�v
Z�Ƹ��ͼn�'�K6��Eg��N=��7�WÂ��d�ߠL���g8�*���ò07���^��p �Mfj2n��o
�?�g�A�y.X��$Nw��sT��:G����җ�*j.�@�ԱMW�����u_}׵�:�k5�-��n��/%�T���$��;Bv0� O�|��5�x��F��+ܫ����C�  |������JS���]��)���3Nj����&��iO��}'��,���z�k:X��&���a�TV��a�:<�
B��A�؜��77u�	{�*���wc�2|�s���E)S���̿��኿r^�l�e��g��ΰ���O���ɩ�%V���������Z��� qrĜxTx��4^�(�	t�|�׽JhL�7� �W�������)�� *�?���Mqq������:CaC��q��f��%�T"��vv�����O,bL�|>�
��{� �
�;�M��,������/|�U������/��@�v����2/S�y�Jr��e6��.�A�9P�*Hr+�j���(`�'�F�FŚ\p��7�o�y +3RԘ�*�Q�������G��*�˪����h�b���	L�V�)ar�d	�ј�3��krX�uq�C36ebV�����?3��NY��^���<�\k�h��T�F�6�F$N����:��m��ߦH��������>���wh�� �&��B]N0�Rw?B,�����tIlv_���5�\��ҫ;��+�v��Ĕ<��܊����Y ʠ\m���	��y�3��k�b��.y7_�Qr�t�G��i���SFN���6�~l-ZTb�� ��=�G����%�
6�93��-)(��?������(�AF���5�l�����Gfh�!	>�G���q�rm� ueS��s��XW�q��+��lH����suڙ^,�cPf�Ԙ�k�R�e�8�Z:�t�g���}3��x�ߖ�G��}e��|z�������]%PZfk�*Rg��n2�O8��m+�/"Г&\�^��i[0ĳ����P=;�s�Qd-�68���i� w˝�Ҍ��h.brw�=��hB�Lͯ-�m�;�U'����gL�{<tm����,z������9��f�Q�Y�.��WI��|����5HͰ��7�Z�)rX�n����vRdɾ����c�Sr�e�K�tAԛ�kjb榈�f,X�f�>����CȈ�I��M�\1f��<����Wi�Á�;�!�B]������(��l���F����/3N�_�#�ٰ"���� /���]�p�l���"f,S�F�a��'�r�6�Ӡ�4���2��F���=��Q��õ6,�?S^<�J'�t��qp�Ra�X�ˆ�i8��7�d�-��zGȰ�/����� G�Dl#��{��N8��
jroTJ��Ӧw7�T��$�roh���:��� #l�F�S�
 �1Z�����|�HP�_�ޥ)��'2&�B����k>�)G7�V��A�)��S��4�ns����B#l]�ctY��0����S�����VKk��9�U:�A2w������!��4�� x�#�L����$kl����A���2B۽��aG���0m��-*I~��ث?���:j�M��i\����B)M�lV��5?t��f��_	��X���Z1}�� ���s����i��>Oj��������XQ��= 	�0��	U��HĎT+���[G��SUF���39͝��x��*-/�Z�1�YL1��x�XT?�|赨|p
��D�QI�H��7�C�Oz�~Bݣ��xJ��)���cIER�鿔��}�R�7��"��{&�6�c0v����C�-�k�#_43gq���\넟U�Ȋ�A.,�l2`�T~���ܘF�We�y�.
�b�jފ(�Z#� w1���K����)NZJD��QT �l)����xB!�6
�(��ׇ��,{�{��0�q���E��5}�7�yWVnZ nX�&�d���F.>mbQ�G�K_G����ؕC�8�9��.��B[�+ l�ߣ�=2��J�o�x91t�g���X�E�](�a�7��|<����"�^c�#���؏6��X��8�Vw	,���Y��#9���}��9/�����i��W{��r�i�c��j�o��t�Z��2�U:���%~T���TM�Rv`���TC��C!�N��/�hٞc}��I���^��t��i���pE1����J�ţ\d��^ʤ�4�P�w�	�Fb�k�A��VC@�q?6�Lԙ�j���)��;F�:�?=>e��F���� .�b�"�
։D��Ca�H!�[�@�~4�����V=]x�t�#����-T� �0����/���$>�{U 
�E<=���Y�f�=��z{���������B���d�Y.�軿w�%�ǅ���2��To�B����e����ђ����q�Z0� er�,���\�ݕ�Ń�w	pk��Q�k��Ӈ�?%/�ci^�I������u��G���m���n�|�9���T��T�;��ka�8���� {���n ��=���<#��VKٚC4�(�.���e�����[%�1pc���/�zH�j���~����c��u�j~cB�=W�|}�cX?[V�!�ΝPȜTU�����
"�w���߼9,�v���2��j��Ɩ媔��A��b߃_���;*���`���T7���O�ȸ�Jj�=3 ��V�<6�Z�QO�꒨m�S����E�����-������Ó%���Yw��l��4e���H�g�X��/v3f!
����=�z_0Q@pWTJԏiR�T�`�_@���q1�N���f�W?!Y���hǁ����'��1�G�j��U4�W}0��L���w�P�z
�!f0̌��K·�
����d�)�&h�k�)>���.n�����ZD��+~�|��{G8��Yb��mg�S1l4��l��?n(�������D��V-�V�a΃Z1�E�U\/K[e�=h�h$fdIap��ײ��0a�a�P5�>V�� a"���}7p��ܪ�����]�#�(E/b�`��Ip�_��ʗX)�M�)��+~�x�uL7z#(����l"�W��.��Ĵ��)ɒ�M��Xx�B3(�$��S��rQ���E)6w��:?V.
���D}�6�N�B��מk�؞�1�aά��*�����Q�I�i���KU֩	�{�QF�+��/b�&=A����l3Y���><Sqn��꽅��UޚI��/I��u�\t��{���}X����٭S��<�;3���`�B
1��55��[�:\CObr_����Z.�u�4:)�ڼ(�d^W/HM�N���3<�F��8%���79_Ru����b0�.t�j��T������tˍ���~���Mx&�L��d%�=��D�DK���n8�gE���8�&�Z�K���Ă��Ct����q45{��E8��1�U��wQu���� ��n�{C%��R�����oz�Qv�^�o�/�n�rΰ�G�E��qNpr��Lk��A��w%B�l4�������eSh�uGz�2��X��D�}ci�u
�Ǣ����M�c�Q�i�#(��_}�F�	ױgC{zz���S�C�~��ٍ�����i%?�������M`�냫`�g���-n)�����Ȫx,��ɫBX-I~v01Wc���V�-��{:C���7���Q_^Ty�W���~%� L�=�j%I(�`�h��~�B��v�Z�KK�դ0�y��\�t7�������)!bjk�p&r��g��������fV1e�6�ܥI���p�qX��^�5N96���c}#TD�:|�.�M0�)�?�����Uc�M*@0 �5�G�͍�0WP�9���f�� ��9�T���L��̈�y���}halFwa�-��?8É��)�v��I�RY�o��=�!\^�4���������;A�:�c�j
�v�;�J�T|���x1�V�X�Ey�򠈋[Ȫ�����qt�]�����+��;��/��FF�Q�9X�ھ�y��9�ŴC�"�)�wwC��R�����)����R���U^��Ie�7�.�]6�W(���`�A�wt,��i�&�G(�z�ܒBn�e�?,yZ=�K�Q�>x.���<��.$D�Ф?�)����.�yuش��;�eg�*�\�Œ�B.��L)�'bx,{|��:�IK���&���zYx��<��@�%�3�E����j47Z�W�����w������-թIVmR+�N�b^�>�������N�d�*�T�uBz�!�/��j�N1s�Le�0}����U����QS�޶�@lA��Ɏ���sň���0�E�d��A��L�b�D��G��%���w(1O��3l΁5�gT$&P�4�J�g衷=u�/��.W=�D�˹��*"oSB��C�_l��n���8^��g!@���������m ��J�]������rc1�z�ܔ�d�ࢇ�7B�~�nCW`!�F-��pPٸ�c`K	0?��Sү��.D�I'�^�q��;�A�mT�E�}��#>6����@���6��`���!�
2kdn�hC� O�P�W��M�,��L�+��(P[�bs,J���1M#S,cg�D�J��f_<��蘠�W�G�H�U��2�'IБ�+�n�ֶM.ұ����tR�-ˌ%�e-MQ�A�/��T6�y�CI�'Q�@ۮٗ{��!-���ƺ��,5�c;�ԝ���ۅ��+����=�<�K�t�w"a��o��DV��0�.��P��^��(MA9�7��ɓkk��Z�p�����[=�;P����AZV(�ҋH3�e��6 I�A�[���HԲ��5��:E��<U��h$R.�Y���x����x�=W�t�D?����&�zN�!��	���4�\�Q�k�%_���J(oF)�~���1X������R��v�̯~}*��f'_+D()&�`�$e]�SUL��߄U|�M4<%3/��j�\�xk
�=��3H /C'ǝ����������<�VGK��+�W{J�}%�"������9��A�Hu�L�"���I�Ýk�r̊��}�:;#���x"̋�>RdL���ˡ�U���7�}���ߩw�A�����c�!o�ɠĪ7��C��� cmJ�Wb��H�^�%9w�7!�I�R�K��Z ;���󷀔�]1]ohR���?8r��`�}�M��~�ZK(r���ޙ��h��T�gʆ���Z(c���}��xL�����
�ж���v���\����SԷ�ό�GF{0�a;ڤ�\�C���p�-����������%J'5�z&�,�kX���	q��������l����p6T��k��aވ.+>a��Տ}�gO��T�]��ŕ�$�-�`��&��A��ms>dة)��8�(@��;�kR��y���4�-v>����-�S	B�pT.��&�B.l�V�k��C�S
|	}4 O��j�'����$Csl�A�	�B�xF��oy��KY(^��� ����*C�~ޢ��P����?�	4k��01c+��Ni�{RMQ��`���$�	����V������gsޛ�QW������l�#.� �R��
I�##��DWM�g!�%}.����E���"��Ӝb2�~{>����Ⱕ}��Ɵ �5>@@�g��|�;"�Z LP��ѐ.E�M�߭yhڅ��7����WO��Z-"v="�αH�Iy3���aM����=?br/�Gce�b�h�S��������]�h�vM�0�������mK�pV	�m:�D损/g��i�I/�r0�6�Ө�Q+�����2gV���H@�-o��{�}7r�6��f�mǎmJ������Kc��ҔH��8Z�0'$���m��j4�K�0�XG�]�F��ka~8�������/�TR�4�˻~�r&&&f|@�9,0%�_֞�r���t���* �[	i�XI�bdė 2Q�`i;�=
t/�TQ��ҡw%�M )t"Of�:�����͈�8��:t%����9�7�?��s	�H�ͅ�Y1�V��;�Z7�H�͔�̉�_Z}�.�&����w �-��H����)�W�(
l��*����h�}@�8�'8v�F^�X ��˳�_��g[ۿ�-����%Ĉ����k����j �O.��x���D�Yx�,Lˮ�X�8����b�`����O*6���#����ES}���M�G�˜x�'�c�x�;��L��
5fy]<\���DR��{£�����¸�}��uĻ/Ϫ���]�a��\P��kn�i���X���)����BV���;�f���a�h�܋>�4Gf���+�r�t�$�7r�������(�����N�C7��t@�m�(�B��=�P�����lKR���<HP���u�B1�*ʧ�	
�jik���NR����
��(�Q�t�g�Oެ����*他U�+�� O��ƺa�%2�Jh-:/H�I���Ej�u\B��ZJ	)�JM�Kᢅ���:	`�Ʉ���e�a�� ��@V��~��B7��LX�o~X��������y����)=z"B�٢�7�֠m����uA�X���1���}?�?�� m�!��_\l�v�ՠ��ڊ+���R���!6�1s/j�Z��j�F����r����s.�o�=��g�0[�(	���D��? �,/����L���M��i��N��S&�s"�Sz�R����6���Z�����L�D�,�0��ܘ��O��*/�YJ���L2�a;T�r>*�o�Q1��[��[O&��T"�y�#��/�S7�fF���S�3T՟�m�e�g� NOJ�q��}\4�:/�=%	z�--���K��L1�cSO�Z��W���˚ي`�Ri�!��w�q���U��l��G��åx�HUI�+b�S�~�*k>�ɩ��LD`�J�h�NQc��D������_AA<Νu�KȈ����s3���6Do���U:�q�_7��;5�V�-��BP�K	�����x��E�g��10Pݟ����6�hǤ���@�t�i����PWM*b�iWPT������H:I8����6��4?���t�Ŵ�N#G-!�\1�d˞�8�$��-�"fAE���e$ �A���Fٌr~�ؿU�u���(eI4�U�8U�9�/���4V�LF��2}"��!in"��K�^�⟁/�3��ߐH>M��ɨjK)�-)Z<"^v�<k�r�L�#�g����m�Z��=��B�"�ʸ#y\�#�����M��ɉ
��,���(���OBąn��Ijm��PBg@����Obp��|k ��Ppnjy �u{��[!@e[�^�^7(�����amJ��+CE(�4�R��!$�n�`q���.�B'椳Jg�7�<���*��FW�s��D���VYlI�f5	2}Oٺz'XM������*�n)!t[�<�v��&3�,N[t�2X�`N����] t.�xp\f��c���D-��❑b<��2�M�5�ٛs۶4AN��4ԇw�D1����N-�T���3�T͑랡	�4$�j��aM�v̋a�g��#U�����}��o���H�go��rs�~��B�䯬n;{/�R�Z�My{{9-���XD�>����䬂X�=��	�"��� u��V��bY��s�����"J��b~�.�c����]�7��*�5{ʍ��۸�6��۞O7Y��������枈o���������D��˽�mED�;�jUm�F���ԁ+�&,�k$=��~���G3����j0)��y%�%�iXE%-�*V���+��Q_�
rN��ڵ Bcw�.��~9t��U�v����p��֓5���e���8��n�6?G�6��Cl���?��mb�5)��y�w�͆dm7��'�%J�Xl�]~�aK�o��K{�j�(����iﱮ���!� 樂�+�y6��]&���dRd���:�8�#A̰�D��_]����Y�!�b_��>_�%�k���Ŧ��Z�OE�|��c�K˫�1!�qy7�9/�Q�
&� ��ͺ._�R��D�������S���h:�����>yſP��{�<��|s[������6͘�N����� a����<��Bt�o	�b{UjAter.B ga���hl�܃|`VɏO	w����OP3$˲�x��57o�(��@�GvZ�oN�����^:�:U9���g�u��lݟ��-B�~�"T|�������O�PHoا�H?����or���Ӌs/�7%�{�)�7O��&i�J�I��[�V����wD��އ�cE0`<a�=�(�9a�&ze��TY���Y��>��OO%��1%�c�$ 	�-�X��[�C2��l�� �]ip�4����D`b5vVk�����~�3���V��2�f�~8�X��N�-��.���S%�Q`^�@��+3���70&��hZ��2��e�?L��c�R����xf'�����Sh ���<��k��;<��r�&�VL�Y������<����pgJ���1�4kX!��ڥ!�Z�~��j�u��U�ʪ���"����~�ߪh���,q��80g(�M�'g�-R�P��2't�]�^!�4G�"�V����@���%��d�ճ�UwF����S@���O�HOV5P����)	�(�F�5��ufn6�T�g��МElƣ돦��MwL���kq{d)u��F�ﬞ�u�
���@�`�_J��'�\�:*s}���K�D��,��G����	�:��
S\	��WEd��	�/<~�3�������+Uf/�,��ǭ��� ���e\�O�%�l���ɤ�k+�ڿ�q��|dY� ���Rv��H@������ ���9�]��?�bj��e�)�⽶S��TM�����g��< ���JD�-��k>��a��M۾	,�P}���pJw��RC\���� x�K��~n�=��+��.n�N��+�-�̒�Du�A�Ǣe�R
��
����ߥ0��~��)�#��8l��� -�X���6d���}����dM���@�3�x��Ax]��+�Q|Y��U�>(ؤ,���� �iPGg��������@�b���(�	�q���G� �di�$�z�
fGuFT�A�'AL.�<���μ1irxu�0� gQ��q�Po�{���;y&1�E�A��)6��sߔ��G����!o
G[��A�2r덷K��������n�-Y�*W/�����h!�W���s���,�KohM�o�%�By'�YA1��q#sI���u��d�OA�6��+�@����-�\û<}���P���n_�Y�y���=��Y�P��"��~?�Y��BYm����O�C���m���x�=���F����؊��Sv�T�&u�����(��"[��W�>�����Δܣ}4!B�e�-.`.�ӓBr�,�O�2t>��ﶪ���z�/��7[���7`~�p����ʰ߃Z�s6�V��Q���vrI�L�!�X ���z����g����a���C��V��#�5�����������!� c�˝KqEP���X�!q3S���� ըi����ܙ����
����%^e���� E��.痳Wv�:�;��m��B;��hWn^-g�;;O�gf]�J@�Rbe
�R�U_A]�y��+�bLfʐo3�
�����������K��x�F�j�	�'�����;�z&S��F���w�Ԭ�C�C �6���Tr��21!�n������ˬ]լ
��=%I9&���'H0�t�4J��>�<Ɏ���I�7�j�����*�G�ʹ
�q(��B�?�{� I�;�'@/�)��$�OϠ����j�$
jT��d�GO���<�{�C�wD�9�ߨ���g@�,��x�E%c�dXTF7VL�I6��.���]��&������n����]��p]v�Hu�b�uM�f�
7Ju���x�,��D*V��4�O&=w����r7r�ʽˍb�@�����C��j���9웕����zX��o�6��/ �{W�ͭv�N�X,Z�Teқ{�M\os�I�Y��E�`h��u�-d��Q<T����g��t��Z\�U��R�л��
�t	��5*ia�˳&�f�w\�w�soE޹��Nl")�I8�����9����fK��0a� ٚ�ql;gߟ�����r���m%��Z2��'<�XOL��I�+m�e]��H��S��`��~~�-2qX�d���A ��o���K\�3&+�T�B5a%O��2��ߠPFD�i܅�r�n��P ,j��om\I+�S׿�7����@[�y�.�?��Z�B�$��Q�?�"���I�|�w%��8+A:Q1�e�
�`��A���c̔�SR"��hk�߫���(Al@�rK[:�\G�ȹ���%������md�|�e����g8 6�3�,���6i�uZU�w��%_۝�3nf���[�I���+�h�,���]�GE��:��_CyN�9,q�Ob�<�)���br6]�l@��Ny��o�{�5Ed8��9ǒ2⢇J�h����-��wA��\-zI�Vq�"���z��n��R0�ck��)�A���`h�C��?��}(�O�MM��j2@�g��0��� �������	g����Ϲ'�o�Ԭ�y�ol"U�4��LL��VMa�']I�Д�<OX�i��73R$+�g.���"��G�^�6���c,�Ӵ���53G:5��.��x���e��YD�{bN��d���Z�T� WU(�_k��0ӛZy�Q����rfѼ���؈�诤�����+�֊�=�vɾ^|��,`S>���П3��*B�=����C�Y"2W��-*����Jeڂ����̙\i����|���BpJ�=<�N�_`�[����g�]��!؆��������Q�J�1�/bs�ud��YAa6 �n/�;�>lq��!��F��6����k��r�������D,E-�͹ŃG�yQ���l������2��������n���Yw���t>�"<�fʪ��W|�����aa'}X�R�����U��/-x&��֒�lCb�М�����p�g�	�u����u))Hv�pRfh������hx<U�Ӽ��w�����2m"z�/P���	���rz��=��+��k{�udi�S�Q7K���Lp�kHh�PN��?�!)n�����-��)u����^���m��ې;i�8�S: cٛH['�3����������c!����>W�GW��.�����؏;5ڗ���4�ʘ�㍊��o ���v���u|�+Ewr����{T4݆M���w^d�5�yV���M�۵-T�7��0rn�>�{)�z�����7�HT,{�[;X'����L����N6����Q�-��6�\j�?X&a�-��/D(�6�F�<��c.��bL(�I�U@=��wn�)�l6��f�..�)u����Ic�Z6�?�6^+��^.���`�Wzf�l����>�р�α�Z���.�x� �2
�nIlh�蠶8�� W)6>�G��P���\��*%F/ܻ��O���)Q}B��1��sf���Rߏ��?���x^�e,d9CiZ#�w�h7���dw^J�F�n��Tj��Ȅ}���R��H�e�XC�`洉� ����"��-��C��tcǀB��z��?m��^�S��b�;�ex���pc[��fn��-���}����Z��X�ś� �	����Mɖ��'��iL[�!kuŀ,-u�з9� � u���h`\A��qM���S}w���dA��q�w|m�(��ώ��'	E,@���qZ��f}��OH����#hb����`7�#��z"b߫�n���*�Qol���a�a�Vc���~���>��Zt+�O􈆻 u�l�\�y$.E�Q{��@}@�����sp��R�H���hb e�hngo�VTg�����J�[7'���'bE�gHX�y<��B| R��o��ȓ]ڹv��?�@5T�[�<.�KҡsCd1ܨ�|�b{�6Q�Cz�b���n()�+x�LD](����5j��8�]�o�37�X��mfl�8�O�AB�S�ȍڭs�ɹt��ȍ�%����l,�%�Δ�4��Q����0��
7\!uk��"3����W�$O��MY$x�BrZ�dr�s Cay�7�}0/+QzN�$�F��"�g�4"��ߝ���u�uT��8�۲�w�i�yIR�H:�e%%�UG}��W���~�l(j`�z�D�q���������^�ϔ.��?�9�Y`��v@(9���]����*���*��?*�G��c�s�
(6���w�@�S�^_WP����P�&;�nt�>�b(������KW���힣�%I+GZ��!X8��g�[�K ��r�Ǯ�c�ÚM�D�[�N}I���%�e��5|���ȼ��memT��\���f ����o����ϋ�	h���i�[Ԩ��*��j�� b����F��3�C?P�Vؒnz���D�ypظ���L6XZ� 6����l&���Y�x����)�|�*�3+h���B�B6����?p��M��f����Z�����!
�� �g$M�l�k_3������=΄��'D>'�v�k���C�_����chh׀D	 SKe;H�O�������ڃE�CN���2\��j�KT/�3&!'@�-��XL_7��4�ˆI��:��A�p��l9
1�u����������\��
{�$k��C�T"	�~?TpI�do��m�gX�nLr�kz���
��[g6�U�p��d�-$ V��,rӌֲպ�>B�G��uQ23�ooo��uwj�K������+^���"�H��d�c�8��l���Áʋ�j���GzYI�J��l�msI�Zf*�s�nS�pz��l3~���?CHoWg}M�Y3T�ޡ��Hv�3k�(ϥ��g0�P��cܒ�Z�����]F��gꇒ�X����#UƁ��A]���_^�Dʚ��]� �.6(�３�7�Y���P}s�]�2��	R �h�?������|�6R�?�,�5cV|L΍�Py�;N�8������JҞгlgQ���P:ϗ�q��������Z|�Q�v-�\�젻p��,xtG�J�n�!���c"��D��h��j�k��e�f�������`M�C.3&"�e�up���{a�d����p�g��!�u|�K�6ͦ�f�]���Y��e�����gO��T�P���b�@��6��_�`rg�	� <tIǳP����;�K�3�o�HA!�0݁�G �\wS�cc�����ر�db �5���������H�8C=�����Y� ��|��Zj�C�q��ӑ@�RK�1B�A������'�⭾��ό�2��9[/��Y��2���3<�h�a���WY��"p5s$�ho*��u�i��$(��(#���E���j��c�w�X��?�^7�3��s:ً�ڮ ��1�w�{����m��2w�?_ɱxc���]�P�� ����:���E�F}�$�u���/cLXک�f����ި	��=XEOk������ �g5�a�.�����@�V��ű�jH&�w�R]Z���.�r���^�M���8ORk��"�7�..��[������H��ьmȼN����#xc�k2�&�.-�P�PX�����|u�5��n�̂�0h�A��������#υR+�BS�~�s��(��g�G�1�,���s�l��(��"�(hw����8ƫY#OS�ވ�]cޜ���hk	=S�r�Z�R��R����4*c�!��Wix�3.����)�&)��2+�=Z���C�����L�3��,l�B�5���WN\��ʴSkW����u��@�]�N�,�eZXY��kf]�Hdz`WK��nI1�/�$72�&d��s�ⅽc'8]�eO�v�}SSR*ż-Q��-�.޸/5OlrYʆ;��<�8���y������C�G'�4�f�7�v�dݡ�'������b�؟ 9��\������b�F����Fm�/a��x��wuHVв�"�W���Ëm,F��S���ݸi�ͼq�)�c%����3�hKU&�'M�� o��o�}�����(]���j������}`�xbq�pv�*=x�q�X�ȵo�S�a/��@D).a��,����ـ�+Ԩh�m_��M�������j�XecY\8�$#X\X�:r��{$O���̇�a���;�}k�D����U�)  {h���:������ל�1��N�zOR+���mb�[����^�bt%a�]_!@{�"-�[��W-�������FJ����K�Y�k^	Ę��"o�W���R�et��#3��^����W��|��V��_�/8�P�ϳ�j!
Z�)Ϣ��C�G��;[fl��>�$�RR]�Fa���9�&�Xe��Ք���$��`{�=�C%���J�+�����+o�
�x�u�DY83�T�����l���`����rL���hHz2�Xv�ؾ�V�\i� (���о ��3_����MY��l�Mؠ� ��ÿ��Km]-�Y�֋�בĔ�{��c��ԧޒJ���;�	�������ҡ%Z>�������c������m$X1�EU���4a�!!@�}��g���Z݉���H�N�Tő�������C2�$8W𪦰s �-��&$Ʋ)�����<�ፘ3u�~>Rp�&H�Vod	Gm��㰒�U"!n�ZZ�e�%Q�=D��e}�e�0MS��Ꝅ�s3b� �� f �6�!ZMpm�Qa�'����LI��eж�i`���r
 �"DNN]�����˧�v[,���Nw�]8���hs�vd���e�ط����u6�Mr� 1�Ͳq�c�0p����X�V�g�A�۪@5YG즇bŒ�)�(��b�N#[�쨆�q��A���1?$�EA�"�3t�\j��Lk��	��7�V�&�StN8A��d>U�X��P�DaX�)In]#)����CƠ Cn&]��u�R�3�8ن�H51I$���`��7�v$��]��.���/����v�^-�z/Y���;p�@�SvY� �l2�e9�<����oZsk.��)���Dd������ZB�<����l�ȃ8y�j}���H�v��n�ʢ|����1�@���m�BG �k��d�sp��@����u`N4��JH�Hi�<r����r.�ߖ�����Qe��S��~W�o�C(L��#C������=�����s���?,��-�a���B�c���t#�s*|�����M�;5hED&˰s�'�1�Hf��= ��,i)�9M�]�L��23��3ALA�汚jhhq������W�-;g�0hȵ��<G6V�o����B���!U<P��{����;N��YbAu�o=3����{@�A>"j��T��= I<�Y��CV�'*a�����5/`@X2*h��L�$p�1}P���$���
���+'�z-	��98���{�]B��o��lT_������ͺY�����!��Q\����-�s21MR���7z	S���z`��"SJ5�o[�k�ŭ,Te;�z�CE�3w�n��]W*���4��.[���.Ě��jI����)�&��$n�s��m����ܐ{<�+��?P��I���о�M���5Ԑr��U8F�+/�go�f�������8jm�y�%�ˠ���תsm7��kM�8t�zDz�d�DO�B�_A{µ<n#�����i�~<�hn��Й2�޹��ԛHa��6�c<�Ֆ��;���,�4��W�4��P��N6�( ��H{�l�y5����&s���:$ &`���c��sh�#4���Ic΁@��jJ�M$ef�f�~e����;��V�?�V���M��n�G��p��,��#H�4�Dg�d�`�ۃ�� ��L���e$Y4	DBH�[�:�Y������p�n)�3Asُi������Ԇ�Mھ��)����'<ڕ랔��2�Z��,��L�!�v����0�
N�cEl�i����A�F�V>���tS����n���c���sS���� �:��gA���*�@MQp�����h}k��}�� 3$HwXn^4m�ﾌ��{2��w��s�#Q��I=�*�@��ѣXJ����/$�䗌��Ov�1����K+	�	>7�[[=P�`w7�C�u��jal�����:�h ���2�fC�����{b1[������)nx
�
���d�	R�,7�'��N����(���U��:JB��U��w�l#�&hm�~��g�][�t���v_���h&Q��rT@�.mW�g�c
����I>r/���d.���E<��%��~ u���mՂ������ز�q�&�1 &��)7 �&��-f�׬�"�3,��"RhO~���Oט-u�ϝ�b�s�g�
��YXP�rHř�G�!�
oW��wd뼅WW`��˞�f�q�W��-y��{�9\������t�/T�_����d2V����38SWQ�Ő�T��(XU�a���������哞e:f<z���h�~� x�D7�����I�;��@�WA�I��y�C���a_�=�V��y�[�U�������{+��J�A@l����j���Kǯ�q�L�o
�ɔ)[��O�	 "�*jB������rg���9�������3# ����ë�T�9z뭥�l�����QU���C��8.���(�̀_|��!�rG����d��t���jS��uj��+'�d��l��-��;��/��� �씘��J��7����7��?��v,�{�ļ�}*ܣ�b0�ʳE^�Gi5���tHm4 �YPAI��E������B���2Z���~�g�����
=�8�#� ����6J��a��2ݼz�r��$�.!�樨��~��Ȼ�%G��tq�6&�£Z�
=Ko��#V�P�oC�	�1:�Q�i4Z�߷�ۼ�vh����iWGm/���t?��dS�Ъ���v�bꌷ���{���+��øο/��hłk��*	K-u�e@����_A]t���ǟp,�z�
y0�_�f��$�w�@W��2�n?|X�ɺ�H��dk�f��ʛ����#nPuH�ŸY��S͎l�Bf~���#v���cj�гU��G+��t)k���nl����6�5����N�g���z���N�V���e\����:l��9��jf,���
��:rT������w2�S؅�^G�3���T����ff(��`ȫE�Q���w��~n�Ho���0�f PB~��>zО�\�8�m���g��`d d$aGɓr9L�iB�
����s����<�|o+�w�ĺ����b i��wn����d�j�/v�Y��uh�=,A~���|��F�K7�l�u�WD�K���Y>�;�>�R��cG2�g���;�,<B�p��l�5�������H2����0����"����n��d�?�R�67:�q������b�(G~�_�O�� a�Xaq�I�ʦU��5��~��l)��`������ʝ�3����|F���[����6W�4�kV+����XC=]�����H��/��Rݏ,Z��H!?���(XSRX*��{;K���ދ�ѭҼ���^B1qi`w��|Kz��m2���k����)z{	���T�̀�F�(��L}IP��qq�zN�]4Yi�����8m֡fQ�w���$����vK9�W;�x �����]9U��K���M��)@E��v��&gɛ��G�@�]����>�`�hV�0�(��'���S����a<W��7./Vh������4z��ﬓ ,!�𘐽E�2�L.��6mX��;gJ建�1�\�Wt��hY��=�K��-�!Z;�{�F�.Bz!��6��,I�ggJ�Y_���VR	�N�ͩo�޺zC��i5Z$}��"�QSޱ�`	�D�U?�a��T�fďl��]eZ~$��cC��z0LgS��
�@��HS'
��r���*�i$T�)��\xQ��=���& ��� �ؤ��L���:3\R����9M����A 8���(1��mw0��W�l��|��wg�/Cۯ��[�ΠAO�:w���1�/�p}���mw����q'K�K!L%��<Z����;]�
:[��W�`|�؄�]�1�\�i�'�A�1��B�Z���{�B��-2N�����^4Npשz��p͛�p�@����>VI��J0�[�J�f�|���	{l���I�q�n���h���y��\w��w��t��[���z�g`W��\bcq�������IF�O�����?��9�ޣb�6��7��'����+BE�?�\-�{
��%/�m��G+�� �A�ڴ�<:���#9�9IOI��[�jb�H�w�����A��w�<mN���r#D_*��cD^���;T��V�/jFc�겈�r�͞�%3��>������U�����?��nJ�����Wʘ`+�B;��z�=0��N�\m|� ��sB?u��ϯ 9E'�iw�FF�%���'q(�޳�m��?q�و�*���pY��<�����
�z� h[,w�F�q�/	���؂��*������dQs�n~|�������RV����kז&��j~� �{"ɝ(�.��2.������J����J��~�xc�h��>&�� �{�*�ޖ�6��<ٿ��G��=�})��
EC�pu�M��9���D4�ᣛhZ~B���21�l�IFNV~�NTC��[��8�v�Ά�=�A��#P�mׄ���J.������;+\�_�����Oo�ՠއ��*(���e�o6�enU�����Y���b��`���\�giW���8v���,Z�T'bg�fІ���ʡo
Q6�+*��]�ð����W'�\�������ώ�Q ZU	m��<a�c{{�_��w�w��w�yMȻ�!�K�l�r%���z��dj
Z=��T��q3Ĵ�Թ���;l�H6��S|^)%��7B&:��5j:cں�Jco��b�����J�UK�g��zg+)�eJ�L��8%���Au�>Y�:�D�;i��ݖ$$���2oز�]���G\s4m"1X��-�t�1:�SR�D�I+��s��������E\x8þCp���.l���z�b0H��*��rd�]͎��M���3y�\pe��e� ՉN��qhW�l�+��\B�U_O��`?z�-A�%�����`�]P�\=����#9j�2�pӎh<l�����Wi@ۡC�9l��t��=��V�|Pz���<7���M��ȭşE�jm)�'�]&����A��^T+�o<`������tD�d1�@��v+Q���ޑʔ�W�z�M�F�����  ���E�W�������xD�L��k9)o. �/�[��{ڶ���j���kT��_g����l�uw��߶e��@�*����d��WM��"(4��S�[�X���:���,B\r죿; x?�#�g���B���#5��Ld�����3�0�,usȰ��x�X�F����)�k(EJd���x���.[~��
=:AY8��� n��Ք�����(N��u���Γ��s�~���֙)	�dh5�~�$��( ��t60+�X?|���9CΐY�ƶ9��d���}	_D�	�Z�r��eVe�I<�B���5-E��i���yL�-���K���ßb,{ۀ�Ҷ;��o�p��ѩ�$p~��,@�������Sä��/�zQ��|�@iG��*/7��`��Kl���o\e�-n-��mGx,���� �Պ	�!�֩��i�|@���l�Οh3u��o��[dڠ������I��n�����ƖWX�φv������;NQHS��H0�t��xY	��\��j
$������@֚� x�"�r?��&�d���nE��E��<PLT�
t�K����~�8��P2wC�����LH�cT����A�o(_��	l�O�(}׭$�H��l��r��HQ�)̩yf�uϿCj:�cCwyX�陸�=��H�@�:ޫ_��K��| �\�?w<��ՙ�7v.��H��%�(�����m�fo����X�[�2y��F֦�K��NlߥsY�'C|4�rumJ����d���j�̒6�P~}wFr����[�KbP�PGjr�?�%Eq?!��rx�?0EΌ�'tw��a��7D�D� �J�+aɠj��̓�c��{�r�f��(Fb���a8
nͺb9e�����^���;����B��dR����ö��0�"u�O�y���Dd���Q�x:n"�s��i:~����m!1�>�@q��6ȤO����u�z`jl�*���jà�Ld[`թn��x~��ź=]��ư�
������i��~m�}�]g�p��k�P��k����?3�q	ɧ�J��d�q0�����A�6��=;�x6.ɦ@�.7]L6���|_�R|�<�7�0�쮫e�W�V���W�B�/�B��며c��i5���O�k�ʩ�:�/��TS
�S���U_0|���N;��t˓�Xͻ��#�]�_;�1�ż��RyG��N�T�js�P�V$^�ǌ�!��~_��<�?ǵ&y�Q��X��Ni_����t��X"nu5� �0�V,�����`�@���L��^�����I��Y�eKOYZ����E�L�	�q���ʈo�炓��'�m�-g, 2L����s���"\�8_!ix�Mxj���;��b��8�K��!࠴"��ƫEA�a���H���A��)�؞"�^�Z����&�}||��9��3)��!s���Qt�\�Q�Y$��������4Y��.ń���s��\b�	~"aJ�|��'}J&��_� N�?�-`��t��3�g�&�9�	9�u�WV�.d�I����A��?VQ5��k8�c"�+@gN�pIT�TFV^c���A%��+rT��Ҷt:S\SH�`�QW��^=��p�)�K_�|����T����K�5���g"mo���R���vE<�h(ż��Ģ�����Sf*
�b��ܬm�T��e:��י��3� �Ǝ4�y	g�Ĭ.O\�j,O�)�����:�������(��U�Y,Ȥ�vwLkv~y��`��:��9AW��ї}�uH��6W��>�<�p���'|q����5�,�"	���"LW�����6݆�r����W��Tre�|�0)�rQH���_+!����l+�&�6	vO�u`бO��jK+.��l��hK��Js[��
K<�,�]���L�9�����ڛX�~ �w!^ؼ��`���T����%R8�:������L���'�/��}i���tB�q�*ɒTk <>T���Sm�+����s���ظ�Y�!Y��Hm�o	'�֩�c�#0���psj|�x�`g顣�KE��'c�Ŋ���r��^l3W���?��G�Z������ִ��%DG!sP���7�����6��PE��	;�p`��9�u�H��y.�8��E�Z�b�q�cB��R_�A���笾q^��o������|{帎�2��v-R�HJ9p덏5Rhǰ����Ƌ��2�?�%�����Bt��-����R�M���+�r%*��oVj��� ��q'�n_$��'nXy�<z~rأ��oX�^�G�!s�a��d���Ȯ؜L��4X��u���04�P�K�T�'��@�B@
�]��ӟ��|6ܫ��:G�w���J��HP�
B��� ����;��~h�E$q�ht��U�|/H;��O>���F
�׍g��>LU�Ѳ9�h42�h���r/�Z���l�O=uݬ�oee�c�B=L	.5��|��j]���w��EՇ�B�/�#����(x��,�-�=�{���mL�6���װ���)�W�f�L*�ʐ��
>D��e,�Z�e%����}�m��i�axⶵ��u�E(}����`)z���=�T )D����� ;�'��B-Hg�K;��=T{�Hftp5o�J�z�u�!�M��ύz� DS��3j�F�����ǵ<��y:^Y�N1R5gY�0��~�	 ���8���<#�<�ƬĐ��@���1�A���O�(1v�>�.�7�?j��w���J��1�=��0G�>/�:/l? Ueծn{�g��l�8yw�Q���!�s�@��^��ͻ�^X�l�K��y�/��@���^rK����I^z���/j�W�L�Dӏ{�?�8��V��pΗ�) �$m�ܾ�"�Ȑ��	^fz���SI�VbA��@��nE��FE�s���K�xo�$��l��7+�o�E�����a~�o�'���|�,T���UT8�2q��7>�tvc\7�o������ih�a��}=��@�l����|��{�M�t�EkS?ф�Q� �3���ù�|�䵛n���E$'^<a�*��:?��-_!��J9�$�Udd�z| !���{is�����Ѧ���L����08Ѣ�皫U����ї�b(�&�[�}po:�a�0��E&0����$�p
r�L�7��0:�XYE���J�L2�d�i�ᶒ��j��V'����w7��[Ƅ��+�~^@[��N1C����Uu�k��,���l�ڨsɐzP�r�3*&?����ΛK-Z��F��`R��V=z.+t������ΣQ���2��U�c�%
��~[��C���y��_����@\�I�GL���%ƹ�g����l���k���
�pt� \�� �f-�>쓴����"M>�<���,%�9�NS��W|uՌ�,1G�P�)bs8�W}P���̑�����k[����mg��ߏ�)��~��`�e���Ox?4fϽ<�=��)�4�p>4�X?'D)���:�/�p��s��|p�;�m{��3u��b��Ot	a�`����r�����f���\%o�a �~֨q]*`�G)�v�*=߃��/O#��tv:��p��>mEXH��q'K\n�c�\Ix\+x�Jcēa^՗�
JU������ � ݵ����x|Y4^8��
�׎�|_�Ѝx������P�5��#�N��.k	؞$�U�Mʞ�� i0;7�w]b!�.¬�$�%"����\[��$kwy���캟R�*�;�ZK}|ڱ���%��S�;85!�)��R:b��*c�G�W�}|�dp\�L}-��Ө��U�6���Tm/��ѮU��Z�cJ��qr1A,n�k�N-%��L��Q:XPM��S��<g��=��Mi C�#��&�����?�	�p��ȍ�l$����|�W���� �>ݼ1_�xP���t��h��)�M�ܹ$��C���U�������B�g��'����.~���P�Ef��esm+(���P	R�>���15݃�u�i1{�ۏ믾�����]����-o�+<���%���4�/��.��ݞ�Tldwc��|W� jG��ۚ��K�3>�Q����bP�?�\p�
�}~��2�����b����5#��8(�q��	q��E7F�oׯ�Rw�9��m��?u�i�%�u:���4�ș h?�fhu�k_�S�(���l�vO$���xt�d�@�!cpn�:K�:�:��ɦT�Uh���/ޘ�<�2u£Z�s��E.
�|�9�Dz��ҷH>egr�q�^so#�9JR�0�+@]��h��"�Ƞ�3����+���ӌcw�|���<�a��j�9��>O�����_$<�|o���㩯S���k�A�A��^&�r�K��]��z5�����[���&��t"rF����S)�$��3[����j^/�I���@]����z:��	�-�h�,O��+�"b�X���@*\[��j��51u�V+��zC��*p8i'�׷WcV<�Y�;on֧vǵ�j�/��ΩI�w�*yћ���A�����遝����p��ǿ�2�.�꧇P����nw���NҴ��T5[��Ĝ�v�M���:��u��ȍ>cU":䧐Sc`�kT��)69	R�T�< �-��X�U������ҵ/��cT��4�:�a)L�	i�+�C�-�)Z� SZ�D�J�y�@�'�Q?'��:����@"u��x���4����XU1	<�D��di-W�4
h�PEϡid�B��q�����Ϙ�aS�!YY�\����:����'�T��)��JX�;�[���[�
{Ӫ�"���kn��� �t���]Y�D���+��F{we��܍�뷓Bg���z�:�h�*��=ht��&���cC
7�,;XlsU�dN�/�i�����}����.��?<�g�ɡ��ub����i �(��͙c�
���`ŋG�U�\�Ծ�3n9�.�����ĒW���Yd@�bU�"��@����5�rc�{�TQv�H*o�<b�{����霾�%���w���Sz�L6a�����Y��Vw�"�O���7$7��G�� �1��A�rͼ��<�&�����=>�?�B#��ܶ���r�ï&i�z)�����ol.: $����'w�i�� ��v��	�j���������S�};���*�s�|�"'6�ӫ��f`{Zv���*}�!ݒ1i�H�d��:8O�a��Jϼ�&'
6n�
!�S� 2z��� B�A�	M<�N5۹�Tˋ�~Ud��bò���S~D*$`.r�nQn�U����ʥ*фxQ�ޛ��]�@�r?OY��_�)�s�=����N�{�Ϗu}f�T٭��c���'��1���z��\��cB��ˏ�t��&����@UR۽4�%]G`,�IA�oe�qn"����	im����~{X'��s��c��j}�����6�Z�9��dcM?"o��<��߃Fq�a�g��눭�?�M')F�A;������Z���q�����e ��D�����5�b'/���@T(��g��I
s��7Rz�%����H�fj�76��H:V��vV[D�w��4_矺��g�q�{ft�U�H�&B
�z��Xy��5��t��imh�$o��]g��/I��sL+������0��u-&uĉV��u,�˂0����iS�G�M����=����:� E����K�Dŵ�M:�"�>p�����x���ڌL��ёG��vЧ�hA^�G�V;cyjJ�Y����v�lI��pc$��r�|=uy�`F�*[�oB������*Uˣ�"W>���*��;d:.̚q� ��$U����l{��@ˏ�Nd���C�.��:8P�=4�R$`�F�%�/���oP����!&�Ъ3j&��Hk\�D�5J�ͭ����V�ݻ߻=�w�[�'T&y�Á��Fp�����uϒC���f�j��ep�St<�~�3�	a�Sj#'!���z��Z~Y+�s�.q�+��t��I��_8y�wG"<}:�.Z���I�`֫�?�D�`m��(��q[J]Ƣ�q�
�)g�`7!�3�܌�9�eT��Z��;����#�A�b����c1k|�ۜ�e��Tm у@��Vi� M�g�̾f��J�[�xQ<�����8���V�y���Sq��h�
��<�b�4o���f՘�	���z�W�k_�?�������F� ��&ҋb�ޱ�Ѹ+�7�
"x�!�٨�f�[0��J��]aa��ӊ[��_�N�a����[D\2��u�� 8Ig-�U0�����X��"CX�X�?4���{J��R����^�A���M�'*}�)cU��-��-�K�ލ�B��J�=��L�����n� t�r��7������K5�w�e����У��6*�����ޞSP�A��H5Mx���i9���i�g��s�b�vʿ��"S���F�C�Oȉ8B��K!��(E� Ss��V�'W���<9�������91��/�Fc�!٨����;��" �����U(a����/�f��Anc2
�ƙK�!I�$��ܒ�84���o�*��F�*O��'�J����3�vl�"3�yv4���/`<f���r�4�
[�ks,�t�g9W��ʩO[W�e=�WI$v!�>:^�������hAa|
M�j��-6x��mI
�8�؁��8��c���&iU��YH�;�_��v�U+��u�7e3"ǮTpV)�x��6f� p���5��!��~0�,�UE,�	���)����V�Q�<}n�
�)�ה��]��.�U�e�/�Q���}�R!�&�n�v J�3�}�#���u'�3 T"��g'3��[ѿعU�� �k(�\X�QC-���by����S�c��L��͞�5`]��&彔�"]7}��*N@*�e�w�"|�'�Mq�*���}�m��5���T#{�e���Y<.On?�wU�,�!芘��}A;���v�ً�^:��33�yE��m�l����԰y
Z��2���R���]'|h�*VM3�'��9��Zw�l�����ؖ��%h�&"��	M7�'�>���}����X�v�s[��R�6�ԑ�K�EiJhExs���u��; ��3K>,.VO-���"�����DT	�E	��f$�`�If�x�����q}l����~�q�x:yv�2���y��ťm����X�+u��G��s�M���N	�;�N��}u��^�rFj�8-���W���/ ��.c��
�P^r���}���r�� ���tح�Rf�b3�;g�c�q"7Qo沂�a��rj5z�����2�0 8��V�?��V+�4G��r}֓U�Wer|Q������/��c�vcvZyC1#�mt辡@�QV�R�\QH&�Ϣ��~:�#�ZG�s[��#�Ү&f8����gǖ��3���
� +R�_����Bݥ�^g��S����s�S�]K��ll�΢ᤔ���D[�]'��"cI���ǥݯ��j�=�]QoyO��� m->�k��@!�{Z��1��v�4��i���#�W�gd�R4��˧����B-8����A��6�"��J�x.����sC��	O�2)O�M�e:r��I/�v�Y�����f�2�)�?"+&$tl���e����M��jܿJ�����ϰ��E�k,��1<�J����)�Ҏ��	U���z��O~æg$Zw�J �����)+,Mg�S�@'���r��Y��D5ҳ<e��&�����nZX������,I�e%f����7$�f���x�&Q�Ig��-���%�\B���6����n;�Sq�Ca����\�O� `����{��^[�P�fu:�������Ͳ��s��������d�۱Մ��y䶹0U��(�|�8��o���9[f��GG|��k���v"[e�G՞�������q��z�8T�X,]�n�c1N	*��/@B�:�V��ɕ�
"X���|s����b�.I�'k�����t�ԧ%�1����R>^>7�q������a��~���!��WS=ƚ�բ��۸��JC�{΋�����Юns�f��_i�Wc�l�Ck}~3��yWL$,8mz�m斋A%�K��Ea���n�v���#��G�u�*���{G�N��r��0g%�a@O0�l���c�z������ڠ�z�og���q�.à7b�3o�	 %}��Q�T�H��lV���K9�j~�#K �V2�xi��H-�����gʄ��g� � #.�=���eQ�����0Z:�y`���|_֭�>JF�T��L�ݟ���⋎�c�?Q-Q�n���>|���n�F�2��[���[L)%G��Ӈ2(�Z�4�i��'�,�N��qHS�*�a���}z!tq�WXdUP�k�ˇ?U��$�gߗkA������b�Z�8SUx���|�z��x=�j_r��s֖ؐ�(�!����M�,���s�M��E4����4Q��<�Oɶs��VS-g�s*�K=4��miѫ,(�$`!��|��W�t�m='��t�!�j�~|�jN ����H��{�t��%��nA`E�*���Qu�!����θ�"i��'d�E�Q"bj�%*� 	)k߉0).�J��$�C$����VY�[oѐd8r����rI�?��[q�۰��%��_�.�7$�e1�b������d�X
��%��2������[��H���lc�~VF�1�x��?�Y��v�r�A�^�U�V&�6�]�_v���\�CM� XC�髝f����}�͕��Gk��� ��ElY@xjg>��P ��NQ�58%1^�f×�5�Ҥ��,�MDT{���B�� ܡ�K5��x`v����ݯ�¶�7\�}�K7\���;)������v�pE�+�f��Ub�gB*��+���W ��L�3K��}a�;xDp�^qڌ� �(���m���O���� �������f�PqFM��=����ˊ��
ҳW
�?#C�#=uux�
�1���7����^��G#e�x��4Z�c]��&�����-�R��Ҁ��U�s"���@'$)),Θ��w#c�s�u�o����x |0�ɘ�r_C�ם�!�V��:���.����������V����N�7rn����5C9;�u ���X7u-=s8/��@kd3��e��3!����SCM˶�W����p��Tr�d7�x�����u��#6i�R�p��ԡpY���1l���=�s��c��e<{�L��0��Eh	~a�+n���jS���~��c���y���.���o�;�LT��+�NM��T�b?�a�R�f��B^�3�R�L|�c� �1��P���C1��M�y`�V���Mϒ:��Y�}��8�!�@�J���?1�P����gK�O�
�-|�"��8U��&����FQ^�Qokv��i$�Z3O0��/������lw�r���6����[�b����Z����n�5mqJ����V>$�}
���'>�I�|�v�_�
	��p��/'�N��)�YŬ֡v1���?����3�^q�x�0���J���|G�ֱ�rc�d�B!�M����Ě�M����U�8�e��<�"֮���m��M�$k��Q�8���m圀������
���`�%*�^4i@���1m�a\���\�}r2��ZPد�2�X���̚(%��mP�f4Qq��K��j[���[JtLa���E?��PZ�[J��%I���&�f���ڏ�B�j�����4I�jS�����~k��Q��Lz}#�(�\&���曕��&����l{'Q�r��q�ypL�s�!�DW;K$Hu��wEs�5\�H�R�:��m4�a��.G����UCz����M��i5�O����� Xpt�]���q�����Tˇ���e��s�QIO�&�˽S����2[��H�Ꮾ���#�Ζ�6��c;�Q���׭/Cc�l��=`dL�{M����P	��1EN�Q�{�E*���5������(��+҉x����C��0�ͬ�8�=�4���P������@��}**:k6��ý�͙��Hs����Y���g�8C40�|����[����gu֧ҶLA_,7�a�'������1�ٸɒ�:��݌�F2{p7��D@J�yA�.BΘ����>z-�,��P���"��W��-� ^+�/����D

�a!m6:x��&�����:�lE�yuG"�c#�R�2G��y"���{���d���z?���Iu�7�Ȥ�l�����b+�+��K�@!��<�v��q��GB��*s9�!��\��/�8sX�?�6GT�xyF���^�����ީ7�����q��P������,�k��0
#o��$JD��lmf%���'��k���B�4'�)O�s\)�!Ө4ڔ��y�ضnI>\����}s#�z_�}�w��x.�"1_U�y�J�'�R�T{�آ	�F3���G�t��\9���U���J�u�v$-ce؏ѫb/k� ���n�.���9�[�����<Joy���ј�wy�-�.y,r�ؠ��?��nr�eV��'�h�:�\�8�u�6�u�I�\;���{,����"n�}�n= )���C���J�ޡ8���.���n<��aT�/[²�%%���Ilj_��0's�"���И R�L^0�;B,����|R{�6jty��fp�1�B��L����O5���&�3���/� 3WY���t�˝?��+U��k�L ��bf�"nc�W��lfu
�=�vq���7��t�L�7X��uf�&�$�lE����叆�A���VSЗ�����Z���(<|a]^��9�85_��0.�LN%x��;k�R{�O�߆�P@���u�'�`#;y����a�Tn�P#x����4�b�	}�;<fzȠ�4'h�H��3�<�4�7E�`?��&�o�,
>��<�욊V��N�l�4�2����[;�G�ߍ�&�(85��ן`W��j.�ѿs%������}�8w'"1��5Ի��E�_ȚJwͱ����**���5LjR^xb��I�MXV<z��T��y��[�[���z�(��1�6,��ы�k��۽;-RK<����M\K�k������Dm��Se�R��w
��[��(�����y��e�:!M��F�>(^����Tr��_��\��@l�
ҥ5R�R�8��mJ��b#�P��qxN�GԴ�簉�Y�}��*�_E�6�
����V� �\BZ�rਦ W^�z�kb~������;&�T�	I��WA)�G�e=��_�*��!A���[U��W^�^7�G���J�"VA�cC��(��+;� ��]�P#c����k)��)��Y0I��l[G���B8����<H&v��K�$����_��,1��w���?`vP�XB�h6�/b�-�aq�����s�����>��O�������cÛu�(Ï��d�Uլ��!�.xu�����<u���s���A����� ��r�h����y�r%#�B* A�$w��_FZ�(:�É��{�ô&��y��?�~Lg n�uU�8��<q�l��%Wݷ��AƖCOCBe3�!��,dD2{�ȑK�:���ɿ��#�����pӅ���[�Vf���z�Z���W`н�58�S�`�:*>��<��AyK�b��I��C`��.ݝ�ua�֜RE�j){N����Z�9v	��ͲV�C��D�V�N9�̏��_��>fim��8��Q��A$TNE���h5��8��Dx<x��3���|8xZ%���Hm7�9��xyDeZ��\�AG%�u�е�w���e��%��|��`�Ҋt��n�"�w;^��is��L�G���M�>��SNoV&iA����J�L�N���A��ǯ�����q��*�*�-���$�/�;�TJ�K�X�:=��0`��Qґ��=ɓK�G�H��i��א0X���wY$Ď�
�� �S>M�@ٕ�NP,�xx&���My��Q��X	%���F�{ɢ�Y�VA�9>5�:��+R�6i/�[!MYq�����4�\T봰�祆s3i���Z���ep޻�?Ё ��	����݁����:K:9�������r�1���\�+BPJ�qL f�2y�G1s<�8�tnN�}u;MdM{;'�:C2*0R�^�sX(����L{�7�97�F�Lwd����P���7�ŕOxNL���Z7����YѬ0���Q}q#�ezz��o'B�aKe���
3�=q�́�t��m1�ܤ�H���:�ݙ�6j�H[L�*��6��{:��ԍ�
�#��QM�`fmByq��Z�� 7�� ��_W;���Y�li�?^S�ILm�dY�W	��� a��/�0�/�����fJ�~HMQγW��2��˜�����y�Xu�ʔ�xW����į�'�ʚQ�7�
���vfuZ�~H�կO�p^B����u�Po��@4��fc�,;�l+d1v�� �\�㕇3�2�����F��}��� zn��读?R��}��y\Or6�KZO�̶̯��`F�����_v�~ct�U��B3?H
��Ν�j!�v�ڃA~h+�)����-�me����}�;@({땣�����q>�|f�9[��\�2?V�ڒP���ڳw�!̜k��'��b�<�VM"�+\eQa�3�F��ne]��mm�6���f�"��n!<�O�C���M�����Xƿ�١��,-�������xs�"U�*KH�Cy��n� ռ&G�;�����D��V2Q��D�mF � ��"�=m��!⹦�UzI�����e?))���ۘ�Vmf[�k�:��i�����V��6�j�ɚ��t�*l�l�K�j0��y�7�}<}=R��5�#�#]��O�`IbD������̗c�= r�ώi����`5Įf��W�tp-����iW��s�'��6�	��9�}�l5!�vtF��"�ݸK��K9V�� �&N�c��(I��?z��K�ȃ-��.�)]eF\�+-���<6�0���FLT)����o�fF��9$.~���]b�DUK���p}/��&0{���~��25��m�u��U�o����ہ�?m����'���2��ŧ�(�ՠL
jN2�ݷ�:��n��r�:"!��'Je�z%��i(�
�Q+\��S�^;sA�kƒOp��'?X~{�	4|��F�c�g��ʂ@�巪oO�y-�[+Y ؾ��W����]����<\���J����!u'��fx�[.")���;ҧAL�3"΂����i'�)�;��p�b#?����L�����+��u�/�y(�V�ݓ92��yK��3D��I�+?ݠQ�a[@�A��ZL1a�.UӶ#k�)!T�AGIм�N���s�L���/�x7od������oUd��7$Ĳ�����G����FL�u��� թ�V�w"c<.������
�<J�$���ߓ��)v��K�Q�}��<���oʾh���ft�U��I�&��L ���F2��6c��c�Tѝlŭ�sVU��$\~�MT�n5(@��3�M�jd�}�M }Ҕ����),�ʠ)^EX��o�"9�^zpZj7m+��C�O��[���[�ӿ%��A���~�(o+v
��KoNO6)��fR�8y?��^ҥ��V����$�p�U�F�� \�~9M�j�u�$'����14�Ab�,-��Ң�dk���k�:ԮH�w��{��d��� �>B�o����_z>�oَ<��J�υD �q����b�����J��oO�GZ��;�|@���8��5�As^�C|ަC9���Hل7=e�[��,�BN&Z0r\�}��:�mlo>8P���kw����t��<��!CX���[
v�������R�e�f�����:�u]4j���:��K����in�\Q����x4�jI&2��i�����TQxW�3yÏ.���G���ǢMu�<���5<WCE���n��WA��)ɚڋRJsӭ<���Ϧ�}�D�E�m��&��ʹ(F�6�>�hY�ꗖ��p&y*]�?]��>�����Z~C�3|��	c�i��_�,տs�_�&��@y�I�Q��m4�j�[=���dC?��Oo׬/3�ѡ�n�t2)>x=��R��Bo�y}K*��_��&f����=�T־���
H� ����2S�2��}����"�
p��+=p6��)vT�8�w �O�����%�i��g����A���;f��QQ������q�h��b��$�!������*3��;��0��v��F4�������:5/�0�&�Y�x�v���i椩Q� B'PA� �ݟ<$�`�����$S��61UON�䍲V�"�­�F~��|r=G�C�ZK�:�S�a�S��*e��w'a��o0�Q�+
���P�e~H�'�)E�[�+���/�B���T�C�P�) �()���o�T0�B�"�"�~=�ԙ�rk	�s难��@�Y�z��V]�*C�m~���P�o����וLt(OY�g�7v����F���^81�o+߯��;���;z:�9���N�-T���}aT���~F�Y�B�V���_C LY�P*oPC#��Q�G�N�陑R%1\/9P@
�	�Ea�jeI��.�	1f����T%��GK�( B�f�ߵ��E���C��FGbA7i�����T�yX�٥6>��������ZƉY���USR���UΖ������3j!�&�	LX��ل����b��ц g@7�����v�]-���9Z�SO��񥊒(�_[�+��d4d��Џg?�*7O�Z�<r$HUF�P=�v��b��%@V��	LaJ��s��~�Z�i+�W�F���e��e�w����f��m�D'��̢�Wjf��s�^'Wy2J�ohj6\�8k��hy[�y�� �L����([$_՗`�GVБ�����9C��ݳ����TV�����me�̼�����!�G"��`M\^�3�L�T�^N�ܢS��-`>Xm�sY��!s��f_�T��f�bI.�r{'yM��3U\�A���[����ĵ:G!a��*�K4���C�ȇ:l&^%m��i�_�u�;���;&��yLT���c������z �$ħ�G��$�/BH4�᭴:�5P������E��Ѓ>~8�����Q	Kqm
�z�]#]Dp��-�3$�+L:18b��~���'��HGKP˳�u���Xu޴YK�/0�NF�:ٜ7L�wk���X�8��):L+V���=�c(03� �g�n�/��ng�<�K�����@Z?h���I�7-��#��)cs�߭��S�R^{.�1Z���
}jsI�?��!T���34��
bdo}����m�*�"��h��Y֐a�n��$��f�Kΰ�C�I���v���%|�o�Z�]������M�QX�X/���\�
�x����օ�7�BeT�J�K���T���]�2Vh�k-��gf��Ԉ��&9r����d��3̛��]�����)%�4��"$P�@�K?%�8zL��}������I��%�Jc�0�JnM�PE"�b2���fx���p�1��n�+Ŋ��=��wd���>*����é��Է���0d�<0��޿.~ɽ)֐y#�)uh�@L��#��fkk)��bp��@�Y��T���欣jgfZooܢe�FIz���,�謬%�&�:-�W����6ߎ��6"C[���*�c�Z�y������a����v[}ɧ�3�׾/+B�#Q�0�ہ1?�����@�3%qC�,�{#�-f�pXUH`HAM�#=��iM������bHD��eSԆ�S���.�W:�q�PI���m�_h� �����ʵ�����Ӡ��Դ�d�Af|�>���>4���w����*��9��Y�s�ƕ+Ec$�v$1��dce2��8�)t]7�%�z j\5 	?�Ϩw$wn�@�V���A�A�Z8]���%^�Ё�U�Cm����a.e�3����'�|z���R)��ar��2���Pk��N�q|��/x&�j5��V�Q�� �q���;YGe�d~��4������[���n��rz5����P\/װ��~�9`㛌�ss3���2$���y����c��(����@1 ��ErW�I���8O���#tY7'wp���M�!B�$��W#l`� ��.�_O��O��sR ��'Ђ�GS�hTR�o&�O,j�s�0����H�a�W(夰����l����>BҔ�Ss�Ļ��>
����p�GZG~�n�h^sn��m�+~�Kݨ��\?���?*3��ZS�]�m^E�46F���y�_@f%L�0�L�6���?���ي2X����S�o����o����H�Ǐ3:��,���>?�O%.2$ ���&��ӦXl��Fl���1��Z�j����N�^<� l�O��`��״�*c��3�y����h�,��C��:��L&)�"]+L���)��^��č&Js�-���y��Z���R'�}�iy�	��:�}֣j=`���Ʉ�W:��W��'����{�L�n����;0{�8tV�.FMX5ć�Hs��9��fW�Z��I"i0��nyY�txC��(��Nt�qb�Q�O_~>-:�s��V1�m����ZSŬ:F��$��5���d�M�0��h�\�_�N�Zc6��KQ:����:r/����Q��`����h��v����5�G����W�w�@WK��I��( � ��)J)�Dg`�E�l�VIW~+��O)���,GZ/މ�m���ߩc`
�Po�fwn�S�=4�%S`�ޖShU���<�(d<i���.Y�|�)�G�0���(B�w�`=�O��	5w�� �7+6�F)D�٫��!��5S���lc�.g(S[�����{��DZ��M@,��K���H�r+~��ԧY��@����4��z1�r2�nƀW2s�m�����A������0Pv�E�o:�Ç�����>� u�
�*��5�����5���\��܋D{WJ>�ؒNP%��d)���nč�<��5Q����G�t�ʏy9&cJ.@��+�85�Z'��9z�Q$�P2��-�`�F��Q�`u#783�uH�d��`��[8O����!P��M�,��ܽ����O�?ȳA�.	>�N����K��6;f���F\��T���cR)~�q�ȩ��#�͕�@���fD�翨͟�F L	���蔳n��x���p��E�ǫz�qv�Ǡ7 ����/E�Z���NSX3@��}H�AF�|e��I��R�·5��y�>�#-j�B}O�	��A[�Wd �dru��@����*�L�\v~(`|�ѩc��f;.�i�f��I��T���ZXH��{#J���,:�����[U\S P�Ul	+Qw�99�z�g�%�A�����|�A��x�5d2}�l�����͂.�pv���*�=d-1O����[/�[�,G�%�S�l����G�h!���(I��o|���o ;���^�X3K<��9%�8[��(3�ݐ3�
��9�,�z��9��<I�D��YԣM<G�̊�~?9��Sn�FVt�_'�ܧ��f���(~�fHXr椵�-��)�b�;�	a�ͥ=��!�ye��1�wk����nl\�C<6��|�[D2AD�"���m�����s�@h��� 
Pq�g;1L�~I��@��3���$g��U����;Gv���k����jN�r��=+���⸅��}����Y�E���0Y&[�tKZ�.F��>u�`{*zԩ68N8p�������i9ҽ��W%cK�Jn�)�� j�s*A�`n��a*5���&����0m�e<)pI�j�0�A��3ׇ�˪��σ?fZ��C�ak��b�z�!�� ����A�W`�F;�N����ZC���ߗ�q��p����s���/�e������&�my���B�=��y���M����I��E�[�F�B ,I��Ħ��-�B5�,4����Ky������y+�:ߤ��K@�)��d/.m9��X��V97q���pn��Q�.Iv�IEW�ՙ�Ѹ,3��V�`�8�g̀A�i�֑��w�W'O�m�k���} ��3��&K�v��kx�s��<:g}'�����]�#�RUW|A�bCmc���Ӫ����A6){ռ�O���-c�3��y����퀶>g�!�L�饇M������C���1#[���=<Ց��E+�'y/��+�A0�@�p��^�9$	A�����,�������-Y�w=���"��$�<:�x���.�v��G3J�/R���;7��/	)��0^}z0������)���0�r��g�x�q�%�9x�$�
o�ͨB���V� ��j��@%1�`�~�+	4 md`I���g/J����6�b���Q����F���%���h��?�����ߌ��i���0t+^�\ц���G	��q1Y?s�T��W���\�C�3x�u�e�m���~o�t�#}�m����ʪ�<�� �ǉP�"����'��H-��ӛ��/a�N^�$�%v����f����Z��`��KonfפŊq$rX��1��aU,}�D�@��95-0V�� a+�c�@��4��!�+u`��)duX���An;�2�����׶L)�	���x��8�p4�OB(z�㥁���C�pTe�`t��v�e�YF�˞=B����|��
�4��*l�*�Qu�zO|NO1����T�� ��p0^H�x�C-Y=�
���%��["��h�`�1�Z�^S�a�7_���-�;c��"qG�M!��5[e��MN������90g(����s
օ.��LTMWZ[��uє"�_�eM��L�t�x�R��e��l`�����4ǹ�y�0���$��N���v�|d�z,�;L�jeL���-���W�{��	�"{4���ZA��� u�_.IxS������Y�B���T{��A����-t�hD��mВ��"j���$N��?���<��7��^�(7�ˑ��`yb��䋔��A&
T���Pl�R��z���1���������%;�k�r��
-]�&��`���*@��
�o��� � �%����H�╖���\�.'�w��*��!�dX�i�)�D��N���z���h���#J,	��H��Gm)P��(��{����[��&ne�a���&���x{���G3X�_B��-6yt��2A� /cu�R��o1�x4en�c��-��ޠ������r��~��#z�	�0z@r>ډ7�G����и�sZ +M�
��x7C(,&��qOm�O���|r��Q���M�	7��������O�.�t��X���4����'���So�<��Z@��D#��D��L�|�1�3��qde;�Tp�*>�� ʋ����u�<�	N�)�����r0�7��}f�9fh��+$��G�	�CgOg�iy��i��:ħ�1�f�r7<��y�(<r�Wδ�U^QOBWV��v���<TH��%�I7�uEό0tTFeO88D�0kD��|zϵ�Ɋ�_I�( �+��>ln��Dc����3�Z��4^��I8�kUqսJ	�-�ڟkY��#Ao�3�XͽF`n��?0mE=0�{�X�Gc�B��!7�
�K�z��(�r��5��pgcCկ�TK�����2����E���u���驼�Ȃ=�Sk@7{^��ꁤ3�g��i�V���v���B{����79��T��X�m�>Fj@^s�нc0"d ���sol��a+ur>u��j�����{8�s b�J�x�b�!��a�'D3}��1��^�*�CDi-Gc�,�?�E���S�͋� *�EV�ƾ:�ޢ0B�f��QP�7 ����Ns�uڕT�v�&�=��&-���z՞���&�V�q�"+n�Ӥ�׳E�;n���b�͜��2�؅��s#|"�i�i
�!���K�zh�0,�Ӓ���1X�]�����K3�[ �fp9�՘_L�M�Z�2���Gҧ���"=S��/E�`��e��F®��
7_
C�O��d�pL��x��Oq���`�pc�������0�.[�*o)�w��D&��)�������7�}�%�ɼ��,ޢ��CuD����0���g�=���3���̟15�����F���}�:
������R�~~:�M�5��v��o[�R-I�~��:�+�QI�k���-'%F7lṙ��{�`<؁�h>�[cN�����<�?{��q*I(����aB�Jꅖr�sڲ��ڽ��4I��x����1��$��S7��_PX�L%��z�W�D#��3����A�*%I>�O�d�#UZ�&�?űKA�XD=.�b��]��,1DV�їL;;��w�O4ב&��dLax����Zf�啰��!�Q����ٓ/ʭ}�D��P��C��5 ;E'i;�8��Z�e����Ԧ�sa͌�+-�]�rU\�fr���e+����7��4�<�B-�l�&$8hҵ����x�S��5�0ң{k��!��%�LC���*����TZ RR�;�*��Fo�@ ��G����غ�NFL��)�?)��vaqi�RQ1u�h|�׼�1��3t�L���f��0�t��`�&��0̎�Ω`:ʘ1�Z�qqsp�G:��&N�k�D�A��Y��Ƭ�`���56�5�1�����W��ߦ�7�,C%z@�����Q�Wn{A!�x4�����lRf��?Z�?����*���)�����y7���أ� #�v�$um��
��
,d���ſXH:kA9�%��NA}��O�%�����
pp�r���׺���K�^e�g�|Q�:|#idp�Htv$�Ҕk:�G���݆���eP��-�o���{OJ�����5�?�hFC��I�TJ�@��v��n�ut9�t�9�3S��ɢ��H���A/��v��˿���sr����Ƭ����ͪ�3Ib��hF�:Q�~����8x�}���K��:���i/M;�ĭ��ţ�B�~Me�'؉����v��+ӌ�l,�+f%��H����+$pRȸ�l�d"n��� �(<���B$�ߍ�o��ݟ��(6W���|�3�b9�3蒧0�퇝��Bb�u�z�Q�8�F�4vR��l�E��3��cX��d�����%�sz!%�k�73Q��PVs<���I�VF�)�)�,��Ǚ�p!L��Ɣ$I�^ �)��5�p���J�vC¸U�*�vW�>���9�H�PU����$�S��җ1�إi���4�p[�L�VE��/%�H����bC�6$
��#]7琈����ʄ�sW��'	��� ���~;$e��9"a�O?���p�.u�*���y�D ��^�w����ot
��3\k,v�;���d�Aq���k��&-""�R�����V��f,p��1���H _e�����6��%��\Z��*M[��BUű�_��1�m�X���'�-�P7!Z��:g��D�\��K��0�:����V@*N0kg'�g���|��.��Z��� ��B��o� OO�*Nǈ%��������I�ч�5�.{]����bћ$��yd%��.9��`���)9G�s�*-�!W�_'=���)�Q���F�h���#i����r#r\$��
�J_fK�+3�2-!Z� �.b�VlD�����2�:�k O�e�w9R��KN�Àz�Cd1�0rC,;N8O�"�q��GM�%L�o�2Ym�?�@��5Cغ-ȯ����(g6�V�1�ON/o��cM,�ؔjL��$vS��-:�����a֯�A �Ya�df	�T,�{Л+I���}��Q7X��f>j.�Rb=H���r�*Ef��iЄGE�je�Lbq�\w�&�>�����7�I¯+�^X��P����. Z��^$ߞLGa���^��?�m>���	!쀋�]��ו*V<m�>�Ҍ3�O��x�IF�� C��:1��_�����	��:f�-���g��^{�)�� !̂�8���6�2X�^7]�Ì���L���磩 ��\��ᄗGEƂ�-�/|9�Ĉy+9�mrȡ�N�_�J�A�:g�L��dd��F�� >d��?�$��l �����{#��׸�_�3lN�z�ԩ�:Gі_�,}�6�`���'���$���H�����n��>�� ����3�^}Z;���<0�ٗB)/�(��c�N�}�m��Z�<ݐP.�:
	��f���_�#��aa�ݔ{��x�Lu��벞_�x����U]���zȣ�ozE�c����cN��1ϭ�CN���<!�;��۠��2"���I��T!7W��떚 0����DK�G��O��]`xY��A�����'z^٨��`ź���s��3���)���[��s��Υ�F��Y��?����z�*�f!�Y��u��i�3�4v:c@8�
{�E-�5Z��ƃ�^ZQ�[� ט2��ʊ`RR�*f���Ey��F_Ό:�x��e�b
���4�\�SӅ�(L�ڀ�>8-��ʆ�����b�_��kA��#��>���6�	y��Sl{�O�n�,ד/|���u�ݨ�𚹿��V�xCռ��ʮ��
˳`�����+ӈ���U�ˏ�0!��	�'���V�gs�+f�[�����La��H}�>�4 ǝ4n1�kW��G[��\�Q��L��/�����"pz��b��T���0c.xx��XL���ʆ-*��Xk����,�z?t��pؐ����q���jkz��I)O�[�'d��k��Y=b�Ǉ��Tx�W�q�F ��F�d8tK���!��X�j���"j#�q�.[�h���ͯ�K��BxsZr�E�����d��I�p���r�����I�o��������dN���8c��4���"�.FQ�����\���Y���/�{iƗ5ȩ�K�+`O�{����z�"���:_À��c[����౺�)[q�3����1W�ϧ ���Z\�g�hU��W�ky���еտ�#�����Cv�5��˗$7ո���?�8�H��z�fށ�fｄ:dϏ�M�@8�@����ܥ"{#�ã	[R
f�8�Cv����QT1"b��ޛ�y}D�g��H��<Dʨ#�{Xg<껫ܴ�U�3��:���f뀣�3��ǎȻ�kczG���BW���K�f��UZn������ȫ��b�,P�ᵁ��vn�}�4���/D5UQ񌲵���&:.�ΗU(���*o3ƶ�	�<�j��t�Q��ڟ�x��,�VYI��Ha�%3��W��C�s����<��	g�	l�ܰ��EST���S��/��v�D��z! �Dk ����@i���Q��:q��(.�w;��Y����a1�� E[���+H@�Sh��=A�E��Vw�+)gp�P���{?]�"@���#W���Ao����3�	B��d�� kAӐՕ����Zn�zi�ټd����� �$l�\�W���ݞ��E`6�n桖�X��� ���A��4����I����ۢ託�	��fҶ����ci����Y�'3�k7q�{��ZQO�ǭ�`�2i*?J�{�h:���o�/�X�sP��	��A����W�"&�z��4��Nfa@b"�Y������ݪF��n�3�z{.~��5g�!
`�d�Y�VG3��:LZ�b�� L�,��5aJ���ɦrϐ}o�/24`���Z��4
��!*�/���5Ǚ�)�d�g�%�1�*_��;�!�Ot��x��d���$���Od���U��Ć��J���@l��
�[�dMGIIn��Bnz6�\;��?5�0
��;�-A�âoB���-x�$������i�!o$a�!7i�K�f疔Nk>����_�����B̔V� ����~_�j����)���@�~�;(E���~�i�|����<៥��f�;�������g}i�@(�-��4}���vX$d���'қ��iȥ�c�B�0r�џB��q����[j1ZH�T���}���nQTi3�t��� iӅM�X��qC��*W�\�}t1�1���vɏ/�+��O=ʨ�x(M��}~��
��W��<#z|��l��)����Z�ᅹs��;49���i]j��� 鬤K�XPƀos��QÞ�[�q?5��ܨ�y�A�}�՗42x�l(�VF#�l:Z��h ?�
6�ǹ/�T���3函���"a�����g�N��c�O�� �j�����\r��Y�zm%y[2&<�DC>y�G��%&�^�RA�����*#�e2�h��+y�J;>���P���v��eܖa�W�q���Ӛ�Z�r
*�t���B���<7.G�����ܻ�ʿT�*�V���e���������<=M3��.#z�ȓ�Ω+pzh�q#F��d�W^��	�E���)g
�E���мC�"�� ,��i���I9�?��IJ��!7�6���)�� �"DW$H6gi��LM�{mU<i�+���]~�C��l>����ĥ���C�db�L���#ɤ�F�eY+j�1֣	fq�
�e�%.�!w�=��8�`�4^��޲Rt�r�[?NWI��������֮]+���m WA"����|M;ʱh��7�Ev8�SkŁ~_ح��$���m� ��]��$�}(�{&�k�^}��p�+���p���,Q0��민e����ۇ�-��]\e�|�j�\nq���VM��y
�t�|�4;�,���?�܄*��b~z_�e���ۤ��G.�o�Wd����JPRt1ͺ`�)6i�{�͏�/
>��&F�lr��9|1�`3+}V�`�_�'5��J�ˮ��`Hy�BX3�)�K	{��nƝ;D�2�WDh���nG�`mo�!T�.9؊���+ϛ}����;t��YY3:��~,h\ԗ����β�G��V^�*��lb��x����د$,N'n���nY�C{�9�QV�I8G���l7B}�����O��� Tp������I%�T~��n�5=i��%�(�؝>��ڏ���������!Mi}ߒ�b��li��v�����I��5��Ħ��O������iao�x��iL�{Gv��u�$��'ȒNS�ԮX�W4ǅ [Ʉoa�ppnV��d�$��o)��˚�H��[G�֒@�A�`�1�5��TB��=���LAIYef=�?XU�����(�����ƣ��t��$�|�IS��*��aq�B_�dyԚ>SE������}x�9]��q]P�G����������8��|�����6������rd�:M����V1�� {���"�u@W�GT�V@�l��9ja��kv��n�d�z�Q��'���iYF��@+U�l�<1�LV~��̝AjQw���?�����S#&ɡ��M��/~��/��麬~��vL�X6&�j���~���CR�J��١��T~��0l�ay�?Ӎ]~:Ձ)0#-:�̶	1�WJ����
�~L��y�֮�;FDo��-���Ξ�Jx�����V���f�퟇&YZ ���U!<�8iTw%h�6D	2�
6��d�f'����r����AL�H���k���^
6\�N��e� y磶�M<֪��"�R)J:|�R$Q��J+��5�؈�6�\\*d������{q���B[�N�n��V;�]�%��<�?��Ǹ���c��Q$�8-UPg��@Ds�"(��?GN����F�.u/*����c4�<D1�#8Di���hz�˱;�Q�b��\#�����ȴ/ĢhU:Dಊ�(aE탥��Y�_`�W��V�����t�^ݥP�*r��K��B�D���U�XhM�>��'R�M�(/V0��h�ϳ�ב$D�u.��K4/) !LD\�j�E��w�g�	yZ�i0�"�kr�r�`�S��������Ҭ.a\^J\��Q��(��(�"V��rh�*�ϼ�y{�\�T�8v+j�e_�zHz��M� "�]�~N���9T�72Fr �р$؏m�hk��o�KZ_*ȩ1���[���	�-Ls�*�^q���O^{l��v�H��r��p}n\�8����`T���Q@���2�����p������Xi�%tpi�~*x`g�J@K$9�q ���F%e߁�NDE��W���9�F�W��g�rk��S�� W����?o������eE2Yn�j.�_a����L����q�a1�z'H��sG�V��H'H��LA䡐}��_�)�B���҈~��?�;m̾����J]�t��i�K������p�Y��5�
q̾+,�ww�����S	�%W�(o�Q;<�v�m��v;�>��Ɨ/.�&�oo2����%2�7�c�cX^�F����{�Y;�4's����By�q��͡ 6�Z��E� ����'&�Ag�7� ]��FJi��`�G����6�`�CO��ޮ=��.���Qk.���Xjh `�ŵ[r-�NI�?Aco]��2S�f���d�;�C3�k�����[���J������!�L"���	��:vo����A ;�-����J�c��1yS�e,C��U��t�s ��5p�*��e�}j�����Ya�xm1���љ풀���XY�T�4RF��}�M�RZ���k���|iè	��>^Ԛɖ���8ْ^h��+����l��T����SW�G������3Q�e������E��'9��r���k K���H��o�`��bd� �(��˝=}�3�H~|z��չ���q��*�G���=����E�W�9�U �m�XS���z,��vJa�|����<�)j�<��0�+=�[�ʭ#�˭�����n1&q�P����o����Z7��G5�����{@���|�'�bï�:!m��I��V���B;�/���L9���Wd���l��9�q�P��>�Cs�f���|��>#�jK�85��	yˣ��XB��H����X+��{
�7�[�����kٓj�}!�?V�o�/�( �$�֤�M�����������9nV��%a6�W
cw�O亏d����W�#�����J� 6m�ǜ�tR�e{6���|���]uM.V��t�ᥞ�w�^�䄃��q&O��^�NPN�):�Ct�wA��a�j�;˗���%A�K�m+�)��s��n�c��ڒ~A��,���Qч�K�����kB<捋*��u�p�;ʮ�^�fJ�þ*a�+{H�+D���&��%���ws�!�/&�̲�f�G� _!��o���^Ķ2�ء�O�^
C"#�+v��/��)��^7TZ'����a�2`׼8�����$q��+�0����u�e=d��&ݠ
�h�Y�wxmu8�;@h���)�^�7-���hW�Z�{a&Y�v�<G!ͭ�K���ߤ��]B�\������΃HG��'���<�8o�eUc{�4x��ӦcK������|���R����rI����ԃ�Y4k����*�0��� ���6�u�p��M��v��J gl+�$Z���0���N[��ܭ��Y?f[�P�m�p;�p:�v�{���\H��R�p�4,�p2�Lx9+�z���`����3F�]SR��u���EľqL�N�Ԃ��7�H [���3�`���f�S��e��_��Ļ��E$���>Cgn�1�3�
F>=f��ME��M�Wc�W'6�ELy��ھ�Bh5�y�Z3Md���GH�M�w?�������	R��s�:�q�˹i�7��9����Rx�	�ڥ�]\x��/�1i[�JoE��A@ӌ�t��H)������%��dtT��I�0Tj�Ŧէݾ��Aj�|��{#<i��u>�I9��t�V �g6�3�D�)�G���C��#�~����J%V&�O�{���7�m���f�|�5�Q�r���}�=o&)ם�HP��rh�K\�<�������֠�ajr��f�����;F�@<*��C�\��5��+�)T-$�z7W @�{�15iέj�6D�imj��|]k4�ǅZ|ˇ�5+�RYmgI��
���A�5X�R���|���կ�h'9��N3%٬�7�D��!~�7���B���m8[X=�E����͜P8e"q�i+b�M�b��~ɠ��ִ�Fn:��`8�)�{�!f[Esi4��FX;P6�.�a�� ��-���ܜ��b�p��ij��̇�W���P����Z@{�T��li���8��z�zV���#�u��ο~�l��I�����2�UQ�z�T�p5~b�a�;��	틯�/��lG�@͹���LʹU�u~u� $?q��&�I�D�V�:�^ �*0������7�*�n��M�h�5�����������#������r�7��JOK&�3r-K�R��_����/�!�����ڦ�-�3����'I��+"����`���|�Hl?�x�BgI_��4ja1����g�V�Lo%��O��o��u�t[�R�F�C^���p�-,�@U���6�!���8d�/\I�Q%o�V�� �z�)��Ь\f���9�����O�VYc
B`08_�ٛ�8�]4i�<�ZF'���ׁ��G�Rt����X��m�%h�^���D�9�d.Ϯ�,)n��M"H6�9_�ąA��_fd�v&ܒǏtC��4Gӷ�`�*7ȏUF֜�r��<���_���.1����J��Q�8y�f�ʙ���<�^��灱'��|B�۽�nB
�G#�F��Ɵ�"��O*�	؟�V*�tO��w���A�]
�-�7���b��I���`J^\�2�TP��W	#˗i�o�z	ٕ{�MD��B㍣��~g|�Z�'�����m���'(�#	=o8��+|!\?%C }f1IҐRe�u���\b7�\���c9+���F�'��Nb��W}V������EƄG��.���DU��X�gB��n���~X��̈no��qv�z�����bH̶���(� �\�(*���NX/��r9�"F���H �v|�Պ
Mܩ����L�������D�<��jf)1�����i�$]��<;V�cB/��ڏ�A{!�s�'uЮ*�䎬N�� �-s(^�E��IՔT��E�P��R�C�Qܒ��mb�W�D�sA|N�׬o�qNs<�,���gD�/1X�v(ˋ���i�y�#&n�M%�Y����g�J^��_�d �s�\����u�����#IӐ�`��y�<�=���Y��=�=�TZ���Xj�Jyf�jzݡ�زo9E�����&�s=���7��=� �hNA6OD�P(�~Ͱ-fk���gv4;�Nw�[�`G̴�N
�Yu����&��W�S)��@v�[MCH3Z�X�p����W�x.+�̚�<M ��e�膧G�5GC�+�}TŤ�KE|0-���r���i�����Uה�����|�7ɨ�/��Ok[�=����A��P�YU�BVy^y��2��dB-Bk���&ZT>-;�(��B{��g@�����\I_Xn��B?�Idd�M� ��X{s.�a�:�� �gD&Mp�Aԛ�pt���T����[��ʺ:�ß�S��e$�$c#1q �Q�a�!�AT�u��%_le6�B%�6c҄l|���[�q8JH�CT�h#���1Y}D8�tQ�>T�j�'j΀�����Nt8,�
:�)��.�Mqī� �'�p��C��lk܇�c� ���2���Ї�K�}�h�o{�@��d:R���^xN�ԾJ�Z�e��<�>���f$&��_\A R'�?� 2!�?g�������`wő���Te��QTć��Q<����c+b�S��*6���ii6���q?�9-8+��x\��OhG�@b1����.=z�X�XӞK(~D	X?>)��a �k.~TC�)z�ا~��4����>��"R��i�κ,D�^B�F�M m����h��4�z�\�M	6��	lY����B���p��a��z�+J$̩Ø�l�{E�c��t�(��lq�u�~k
�5�%8u^Y���Iq���c���Tޡ3m��u��6�e��}������]f'޿(�K�I�ϲR��v^i�D��������YT�S��`���V�v|S�_k�t�?�UT0W,L��k��X�4(団�aY�V�o�6尿u�=&"�k)w��̳��튥Fb�:����ϘS�%@�)�Gr����Qƕ>u�~���E帨e�Z䈔������HG��*��p/��b�#MP��3����1,,�#,ƖU|�qǟ�'�a-Ǐ�A���A��4�#:ł�������4�)��	�h�*�'�?�Ѥd*UE���嫐t�[x����ơ�I�F|����|F�[Jgo����UG@*@ۤ1��z��~A���%
�������vu��K	���Ͳ����+D�����/�.�6��F����/_W��8N%��� 5�R�覠z���ؠK�z������ئS)��,ٖ#�l�J-���y<}+H����}FO_5��E�M���h���%ʋĜp;�B�(j����6���l���*��{�Jh{d���FZlw�k���ǚ��ިxΦ���~x���z�wɒ�y�
{7J�Hy��e�YI�S��*<�^ms�i���ް��M�x� ���VOW&z����pZF�V28�y�I��AT��k�-B�H��t/1ؕ�iK����<X��ɐ�\�����v��ʋ��� �%@�Ӵ�sJ��A4���ڞM�!�jړ�5�U����k{��ލך>e�;����b39_#�2��W�v�-��I�?�;��s~�K����D�G�-���Bmv���3<�q11�1N���e$�_ �� v ,��՟��WpL\�@ީhP��P-0D�����Y�.+��c����e��� ��?�/Ł�@^�
�QjH�#f�vA�,
�?�|�O�۠Tl(NajV�D��W��V��Y�PdŸ��_��εC��M��$���MN1��s'�E�&����jӻ�j��X	���>Գz,C�:^Ǯ����9[�af�����:��*�i�oG�88�//���I�d�Z��D-:sH��|p�r�����W�7�������wxH+�:$�%셩l7��2<�JcMӑ���[�����f#�݃hL�L�$�E7�H�Q�'�}4� C)���7̅�&����G���wb ܊���-�W5��^�NJd��$�?e���[fJ� �/0hL�ë8i�r�X�_Y�H��/,�J������k��K1`E��z��5�����	�Ė%*����Y�*wY3e/{$�<�tLt~J\B��jy���e�U0[ߔ�ƹ�8�n�s�I2� 1��m@~�Yj���;0"�SΠ ög�����Y��Ǟ�̜#|��S��E�SO!3���6�N�z�{�lBm8?њճ�鸔r�D�d���w�% %'փ��G�;oY^T������������B�b��-�ˠ@�بY�I8j��Ffl' :����z�B�U������쎟-�j���F֞�N}���B��KVa�MB�����AԘsv,N�I�
[u��z�|��@?�$��1M9I�c��CAI��b�Uv���P@jGz1O?;ER�o��B�	[��,b}=�1����}�$�[��]�4�K���n��eڎjL,A�xV��R
h:w�׬�4ӥ��l��ܠ��rÉ�$���C��MX]����<�e�<��5���tV�#+��yKu����:ά|�U;�I�������WĹT���.�5d�uiM@h�֙����O��f��}���� '��]�w�q�֚J���`�"�0G�"����vzk������`ΤݩM���$7lS_�KN���������e�[��D���2m��~}���J��Z��e�o�a�v����r�j̼p�d3�S�TB�n�%hQ�UGep�qC�����M�X�J*�;�����6�/���J��6	o���ݚ�le���9n���KRi��`�,?�i=o1��m��p��}2���{LD�)�V�^�4J�ZH�=����4�MNS��f6ˢ=�2��݆nW����.�an�7ˏj3?f���
#2�y���1�������%^2eÑ��vk��%�bc,�'2]�ҙ�x���D=Ӏ+I9*���$_#w9�h ]،���Ф�O9ȴ��2���%�#9��Jx�O���ИS�\ �{���<M�eB��4U��'��\�B��,���x�����ŷ	�*>��l�pN�}�do���p�2-����#m��H�?1�x�x'R�t�Yq3X]�Aq�5S�nI��DΎr$�/F{�?l�[�
cF�B��iJ���C��I�.&��c��i�H�w� �S�2�u�P��0JI���SސbY�"j(��:�@�:�Y����>OL0<�����o�u4[�^�T���	
9�ٗj��{ZC:
Ck�������R��Q֕|+V.����~�1�@�_���(��@mD�U[�AU�2�+��ly�c(�/m0jм��I�?��N���y�;{�x���>��X�����?q�f3�i<�@�с�Av<Kt�zB�j����\��0��Aa])�C>]�c^5`����WU͏�d�����;[v��f���J��ˠw&E`^���kC�/)�tL�;7"���������� 엛���t�5���P(|.+���{Q����P�����rO�릋���5S����PoM�x�yJ_C=@�wS�Y4�6���wJdݮ�Ƞ��K
0����s�ΧZ��Q� `K�&�a�������K����#��2X�sU�y�6�$|�e}��c[�@=g%mEn�l�E!M�z�+������G�G��أK��+i�ѠC�G05��?T�pR��~�)�%`}K����w|�V1�#�Fn����>;n�n�[2g�-=u����uJ�̉b��.�� ����Y�ܐ[�>ʏ�6������l`�0�c�B��^3{&xER8�\�yqi&
���f}ĵ�lHEܺT��G��5�;�l�@�%���@4�\����2�[c����e�^�/�s�Lɇ��'􇗶3�-�f{��&��B��Nrč�_��U}Iv'��l/m�LydL0g�6�OQ�'(^\�RWv�����-��=��5�P������L��W/°ކq�$�]5������p��U���Mo�Ѝ���~����=�3�y<
m�w�]^�[Ls��_����%��/,!,=���=����pR����]��6��A�~C��o��	�e��hy��kS�U�;�E���g���4��W�����Y����-=��/�S��#Ո��ٽj�	Z��*�3�(�����#����4�
\;u�@#?/6h|�x[5��
S�w6>��L�	�<���c��UڂXcA�<��4�o��rMq�V�e;\a҃|���cV�%{i�e��)�|a� 5�;�@�<|���܏�B��o��oԬ������������K�r߈i��E�_����t��22
�#~V5po�������1D�y��'EM(�/�q���yJ�Y�NS��49A#K�Kj�+K�$�/�3�a\�A�]�W4����\q,s9�`�*�3�b�)(��}�����errX�2N8	}��H/���`����d�7
�j�*��3���`�ؕ}��j�=�<}� ʻ'F��M��ޭ��"a x����?SǑ�f��[��udf��r��HC�"e��+�
�6�~��p]05�7�^ ���g��dN޼�
���^;�	����_i��s�<� t�F=��[y�j�m�7��Qq�Y�*"�����r�K��B����HW.=��'Un)ۥy3c�jY-|�9
4� �"y(��.I�ZЭ���?�D�k�K�-ȯ��w<����O�y4k?
{�ח�f(�d�aol���X,Ho
T����:5FW�8�b|�q��=���$k��>g����d�j���Hpř�d'=h�2�v��$�G��c�����g&`Ƀ��V�!F� 	�@�=?����`�A�����;�[�-��IR��|���e%���
zC�>\��&���v(ˌ����A�^^[�@
Y�c���J HO��^n���v��.����Ù��[[�,}ͬ|c���K�a鬲0=��H��М.�D	�H�P'N�ٴ�c��{C[�[Ml��>�09�	�sI�OeU� mc���"��݆��+�se�N,aZ]�Σ�0բi8	�������u�`��>3�xO�64���#F�
��P��B�6�;A(�su��l`���3Ğc���!�k�&T}��u�A�y�-O�r�V�?��i�0�i��@;ˣD�p$1���C:�H�a���ăT��f_�=<4sCc��ᢖe�c4�����#$d��Et�5��5�ڄ�p~���@!3w�+R5�,6\�hf����\�C��f��?�t�B՘�u�<�Ԇ�Ml�g%�K���|�+���آ����j�dJ_t��B����[�!@Մ�P�,�ɮ�ޝ5R����4�D��*��5��i��Z�X~�aca�?o�o�:���8<-�xve���j^�Z x�+���r��MU�XȠ��M<��;��������p�����3@П��M]�h��]��Ǒ�ƆP�U��Ԕ�rP�@��q]� �'����/��1�BNF���Ǫ��ǻ��`�A����~��7��y֚�q�2��Q�֣�~�4���gԐ�����F/�h�y5�x�8yٓ��'�OH96p�x��NM�:a5LBt��m	�;��`NE�k�gl�X��kӲ��~��?��հ�1�Hv�6�w1��^$,D�+��4��l��T���raD�'�x��ZxEQ�4�9b]>�m��L���I�'�=@��î�(�ѽ�Ҏs�/rS�N��H��D�uƩ�xF��'\	�i�A���ah���n]�z�0�i�-{�pd���f'*����=7R�x�gQ��ݜ�"������*�}���ۡh��U^��r����Q2�NJM�b�i�f�ƾ�م�e�Y-!B1�r}�P��ٻ���1r��_��z<��7�\;*����|t�8�^���iY�Y��3�+B��ڱ"� ��2	��:jhJK�)/?�*�긒�&�dK�H�ڧ�I��4:�=D��ǈ�f��Y�vN����Kn�t ��f���{�^T���o�ez�UT�q�g@���K����Ы�
�d��Ƭ��!�Y���ŋ>ɇ`t��3Aj�+nan�X���`X�uc�VǴ��S�E*�8&hЈf�^�m<���R�w�f��E�`�~��o��������L��T����5P�Q�v�d����Bn]��͔�A`O�H���{�oΛǀ%{�!<s�g%�7�?<�rL��P�P3G+�h\�;!��7�����F���﮵�jt�\�Ă^պ@U��J�Z�d�"������ G��nȣ�3��_�i�.ڮ�5���*eK�!��}�zD�B�\��}]�B�[��F���E�O^F@>z�=�;?y�3���+h�N��E.d��aB=ԫ�c�m�Ĥ�}�N̟�Y��X�>A�u��J`	�����|$Z���J	�\'[+�jxSÈD��2�����t���Y�0��dg�p.���6�괴J�>����0_H;��?G�+�Ӹ�0Z,�;��NL�6J�~�`y����*�D�a&�-���	���/g� �
�n�kc���4�������=F�`(�i�Î��N�����P�!j��j:�&�`�ⷈR5�"�e�z�_MBg����g�<�����������%��%�}ʵ)Z�#�
Z�����AP ��R�( ��֖��8��x�g�@�gV��7��1g�|1�{pF��XJ�<�	�-�U���^!7�c˞p����X)+y�-�'}���Գ\�]��nRd�]+��G��^W ��>���U�vZc�@�c;"K<U]����ѻ2��<���~`a��GF�f �&��g��C$?� �<s
�9�m̈́�@d��vΚ�h��{�z�Ğ����puN6���d�buq�"��
vaփ^D��䣃<��!�{��_�ߛ6=���q��������X����L�ֳ9����>��*v)W�aYi6��s�m��P���e�Pٶ|3�>>��b�L��e��om���(d\ܞ{X��\$�N���~JqO�;˦�f�}������3`�F��`�x�!'D�	=,Ž\�gD����s�a��/mk�Tào\<��|����1���f����b%:���o��4#�tJT���8qwc��2��,܁M�K��t	[i��V'��^�aĳ�����g�E��U����G�<���cˏ��e��@ۣ� ��rt8|�l'H�={<�<.y]�<j���u�&F������5��EA�������Oo�R^�l��D�������r�t��+��#6�����90%0�U�U#)k���P���޶��lh�Ik��3�e�f���������� ��M�* �T�y���w����+@⼰�	v%+�M	%_��/ډ���ؤ������,n�Ċ��R��.�����1��x8�Ώ����5NT-/�1sA�i��tP.@Nq!����u4Rg���a��B�򰞤�a�Ҙ[N#�c�wA�\��e�u�P'�S���|�C�A���L~�p⮧C�7'�T� ��Gv�j�d��b�o�N�s�Rxl1K�'�U��;�^�W&�����ځ���ȇ�xxe�����c��S��HC"�9@�G����7uK3���06�ٿ�ڮi��bKH���f�� �	hc�EA�"�죛k/@����<1#�!�\dUaVqx^o�86��#v�~�U#	�\5��+-O8 �������Dnќu�	���VTp<���C�=î�x����a��>�ɱ(_^;wSw1���� � P
�P��&�B>{�)DF���=$A���2厤��ǝ��;�/q���#�H\���=���Az�vG���?����I � K+��ђR�W h�4O��O%�^��x76X=Ց@j�H�g&"X�ZT�_V-o;����-��n��GS
�sL��KLd���*��ӗ��YX�Xq����}�I���>���b	�q81�.۝٠�Ų��T����5�k��"��?;Yҝ5)F�~�H!��(�C4/}����&F�}�fa�y���=v����#V�K?�Ʈ��`�������<X?K�c���݋u�Yb��uG��!
�)g�a��Q'𽼢d����7jw!=ȏ���5�pɲ<��bn���#����2Um�Nv��/:����UJ�V��@�VE��K��Bk�&ĕ�2z�V���~�Q��1�z�p#�Zk=1�m�X�ה��!co�k+�6鹝\qY���J���}о.�B�t�D�'d7��;��L͌�m�GvKI�F�
��Y���~��ŏW5�F�{W*��^~b^5�r��ya�![h��d{�2_����$�՝bŴ��9�3�iFip;��n���������U����ǹr�O�K�!���#\�=HXx/ZUt�S�������^�r����#ю(8?�H�N�@�����he�M�;պ�~"Z��Ct����k�5C�7�]�SYg�nm�<�Ű;����ӕ�]���OU�ԫ�S�q7(ϟ+y����^b�C1�쎍�s�sMy(��:A^���`K�P`�ɔ��nn�KH�7�r����B�$�?���l��u���Rޑn=��f ݥK�������1K�K�+W��  �]�,�<�
6�p�]S��Je��i�P�2�(��(\nıP�rb�$j�Մ�A�Od�%):6��8b�J�ΪyB�WK���!��V�O��� �Du��mr�h�Yx� :�[6��i|�3+��%.��2��R�m����iE/����^�ݛ3���a9��%�?�Ś�v&��f�ՈS���3�^7k�,���Z�tRZ�1��"3nIC���=];"���k�b��	�p��d1B��p��ӸC�~CQ����<���ӑ���ܳ$U��CD�>ۮ5�;���o
�h���x�͛��*���B֪��8�~n�"�I��1&aW���J&T'��M=G;�9��p�=]ȿ��ډ�1|���7m��A8��O��N�O��)jn
��u�K�*�NvOS|e�[l������9}�K��o��4PT�Q�����?�b���8�3�%�ln,E~:D��߆�����/M�)�$4�ʋ_�?���:jh��4>��kg���!�k��^7rB�����[֐���*;�
w<|���c�r� J����
��HF\�"#2d�<g�B��Rx�����/�>*�����1���5��2P|X�bLa�PyV�)U�����"-1�4Iz�B����k��P� 28�0f�_d#w�L_�ǹ�G"c�=���p��O
�Û�K2=o�
٘n��ZaЁ�������y�[\ux��V��zhc�Ȇ�Ip�F��	��o����fK^����g^���`oM�Ȅ6\����^�S��2uP�VE|\f3+n��j��0����zl����ߝ��L������$����N9�=�k��fF���9J��d		cc-����ç�h�`��q ?h�Li���U��@��u�nj�cu�X�̹���W���V��q6#�'f�`��
}b��-��9��~���.�q�>�Y$�Yf!����d���dD�D�.�����& otr�0gFQ��rU�ˉl���-��#����#��@K�H����]/!��`���I�)�i�h���\WO�#����9����{�h��O;�H����u��l����^9߫2��<: !�ر�f�=ٮ�f� ��@"k=��KЀ͐ǅ�	��ѽr���Ld.ч��\p�c����(���t��!�?�"�҆������0�$������_��fw&,6[f��A������d�u��킗��Q�-�0:��yj!�|�A�������Y�Ŕ�r[D�~#��`��IL�v��B����l#���s��S�������o"�|;;��&����ۣ�AO �/�>��4 ŉ�п?d5����QK��B�0k�!��n#["M�^�bZ�#�9�O����ڪ�ͣ=7Ƌ~��oW��:�̳����iza��.�����Ȑ�[�������cV��X#�Nd}Kq=��[W��fǸ��(g��Jz�G��M��+/&�"�|�< ��,oBnBۙ��j]�9���zr����"xӧ�����æ^��<D&]�K�����ӫa�A�x�����|M{ѹ���W��
��t7��	"J�ꈊ+�X�f����2�%=���*4��UdD����ax_R�F�2�Rw�Ѩ*Yj+VFT����q m4���DR�'�4>�X�~cm���p���v��7��Ӝ�2l;����:~	�ƺ�/�~��J�[�0{�"V-~��S<�ݣ��m$)��n�a?������:6(�5i��s~�W1�K�"�a���d�3d��'����������i4��=�eｔ�-B��A���;f<n��7��D&�#Cc#�^�ʰ�\�� ߘ����ݦո�x��.��-����v�\<W��3��1�L�,�-s����ػ�K�Bs�h�pȚ����ݼn�Xu�/ L�r�q�����Y��!p���*��K���o0�noJ}��Š��[JYvui��d�)�f��~T-�HQtQ��6M�ϫTw!\� MN��c�ui���޿.�cr� ���S�f
���#�?��dL[؇NmA؅�P��j~N�~��	v_䶦 7�Sw��hừ� �MP�j(�'�&K��3#�48L���ATԔ�,�B���(�0���Lz���7��XA!GYjF�m �]���"II
�D�\�|�&5=p�t
���	��m�2һ��#!`���W��	OI!Mu��:]?�5)w)������O"��hMv��W�����ď�g���
2�Ƿ���.,֬޳�;-�H�\V��uG��l}�W�������3[�����<����Ʉ��.:e]��v�xڋ.�����wJ�Rb�ʢQ3�ۊu�f��~��
�*jA	��_/w{��8 �K���:��W�?l�~KN���"��Ozj�%�S;�6��^0	�vw�iy ��$-��UkI�j��"	�d����o֊x~rvK���'p�()��_&BߵG��BX?_���de��8z㘑�5>�^��ᨋL�}�13?��e��@�>��u+��Ϯ�½e���0�ط�m<.;�؍Ee���C: ޝA�i_/���> ����Q�����p�E�%P��'���c0��X\����hM�&�ᛉ��/C!�.W�aO�a�x,��Ѫ�U���=[e���]�uǬj͊;4ci�R��W�aJv-)��r6>9�i�͸�=�궡WOd�ԾUA�����@�7Ud}1��ߒΖd�`�Q~�z��=Q��hoi�RK��4��8��=�K�x�*���&S�䇅dѳkW7���$�b��̾Bd���,�07�]�k�Ѹ����g��W�7�l�h�T"��@nE�J`‣K�����#�1Q�1h��qX���Iѥ��n�X!���2[��B=7��l\@��^�� �®����m\��8و�);C�)t]�	���'���m�ܻ�&��_њ�)-������)��p$��b�e�,:��5�/�%�����I�C�`��C������gؓ�0��b�rs:y��K%n��sD=N��'�nI�B��C�`�{	N{kf�۬�������u���4����u�8��4��7��*\E�UÂ�gq��Ef|r��5��P�q�4ә�b��1��%Kz���6>��\�HO~�*��ڎ�T�dp�]��7?m��?�AG�ʅ���vpƻ^^��-���8[�J�)�j|P0(�=�N.xB�%��u�<�{�5�۾٭!���q�O):��`���طv����>��*�V*<�}�~r���$Q����p�_G��y~�n�Y���OZj�4C�\h��YZ�������%-�vc �w�A}}[-���|�J��*��v`�0���u����@t�ްm) ������m��ҡ*Z>窅�ꡔxݪ�H ���*µ8��E;ǐL������������Z�n,c��ъt$���^�{9b4�#1D�J��H �Y�_�|>10���r�"��"���0Z-!U1� �5�0��#_��Pv�ƌy�
S��i":����N�V?NC, �����PB��m��Ѕ	m؃�5>3�Z���*J� __�Pq�S&�|�܌�%.T�Z�$2/�5$�Q��[���7ѷFm)��Fl�v^���O��z�`����*	dA�,j���xbE"4id���w��Ёޅ+��J���+$�b�@Z$&���b� 5���6�1V�����V�իM_A��F�A7��6�?k���&����(� �;w���#�F3���nk�����iV��:�g8�����b�QQ����\���o��B�҄рO�A.��������R�����ZgfPz9�J_}g�h�\ݻs��;�1$u�J&�VJJ��.zV\�R
�_U�|���c�V��uq-!��6ԏ�����$O�j|`���pl�^��50E�b��!*�,r�S�l�l�Q9*Ĝܙk�$�g!<_H�Z�H
�ï>�ȯ������
G�P������ʐ/��x�ǳ��v<��6���{��䭱�����Y'r�U>�/o����L>����}��v�`a;|%�H�V�l�������lQ�iU�oͣB�lh�z��^�ׂ7'��`s�yZ}��iMk-�#d�X�Es1���Z0��Ϝ�,\B�����i)��,͔�e��v�#z`S��*�-�5��'�u:�Ө�~��A�,�B����,S�O"����A�m谛�V/]�twG�o�����������c]����%~�LTP�
���h w�4$:����H��h"��6��4JE:���z�	 ������ln��V�z��J�!n�sB.޻)Ѩ��$���~p�.�ʀ��ɖ��R�my�Mg���L��#��C�6�|\����|�2?i�+\6���gV�7�9d~+ߡ����Kᐥ�W�-g�D	�~���<����f�����1�����o���a�$��m><�ۋFKlY���|���ik	����Wֻ_���S�{��F�nx��.o��]Ċc�Q�����]�+0ͬ-�ҭ�{�8_����Q\"���$�@[�5�5���>:F��=3���z~|�u�eEİ̺Ze��oɜ�;R�7�^h��U�5���T��y2��wT+փ�xQM�V��,7�+�QaA$��kB{�U#vW�?�����pM�}BIlb��
:��b�<2C�u?�#��Mg�EQt5=��zʀ�'Nm0j��2ҝ����9��l��.2Ԫ�}���ݼ���Sn$k>]� �"\b���6�/� "»p�C�ͬN�_l��i��%rV�TK^1��[O���V~�4�V�����EX����KT-)�^:�xt����!v� WY>@� �)��W�朇>!�BY�Cy�,_F"�8G��wu�
<cl�m���#�-"kW���6v�l�`��so�L�@7M^%���9aCĕǮ�ƶ0t�4w���ܷ��D��J�rA$ːxIM��Cg**4p<cI��AC�[v�&&�4�!����+�Z����z���۶��$4���ǂ�����éJH�T�?<)I�I-�Z�	�+56_�~y��c��W����Ym%���J�k�W��G��[v�9-�)D��4�f��ZdÐw;��z�i玏��Ze|H��.a��i�������m�4�qġ�W�]�z�&%ws=wV�;��H�<?A���QM�48�g?��:K�t�1E��/r2�Dn���_��8���~���,��c�G?q����L�౭�4��e+� K"饥d$�U��,��o���|k��ْ�6�-�%����4ɶH:s����w:do:�$���0Dj����L�$�H^�#�'Bn��5�$�$�uÌ3�:e=SV��+*��|�{���`ߛ&Bf!�Q���&G��&*��ͥ#���on��(]�U���/��)��џFM����H4�D�ڧ͈�w	^T+�]+~p�e�Wj�L�C��y�&�j�Y
ո�-����ż��{=���C�m�u�*��A��'ĉ����r�M#�5�����Bn��e��� n�'�.���V�(B6^ p��4ކf���g�����"�C��u��t�gU7�:�%Op49�	��<e�>Cy>t�<^@�B. u��m���r�E����Yr^�0V�p����)dx$��eE.(+�\U�p���tr�U b[`�I�ۄ)��C�J�G�]s�hb���z;����`�����t.�=���p��N	 -���]k�Z� ����D'���;�`�d�q�>X��k�i��X�\�D�
AlJ�� ����:��@�珬����̲�-î�<�s��J0��Yf�^�S��~��.B*���P���I9��u�U �uo�&yr�<Vy)��Y�s��N��w�X�a]t�e�>=S�!���X5������I8�E:�S��PY�k�v���&-㎘�2�@����3�ZW��^�ot[��ܛI���AW�S��ԋ���mr�v8�<����ٸ�Y����g
�l9T����#񯬥���0\�����qZ���rE1����_Zqn��Gs[���U����(���V��m���c���"�n=	!IU��cf�p)�
�+i�W��Rϥ~&U��-����M���OX�a׺�t���=V����[���w�ĽN�n�T��+:��m�ͤnu�U&kH�
SB��L*N��;ܾ��/�Nk���
lV�3s��e�#��(��I��!?��|RV�R:�0D!�����Xa=�"~�3y�L�)e�+�bD��sNԩe�(ehA�te&g�<eU�k���t&7z�%s,�e'㏘��O0�*�s��n�b�[��6�:����$!�L���t�?I7���*���D�����~����I�%P����#�Y���Lh�J��Ub����)�1ƁvZ�� �/,�f���Ϭ���5^SG���R� �6��s�/ƁE�+�����vc�2N?&Yf�%�2RD�����Y��[P�嗽+ﻏK�rȼ��q9!S ���-��#���ڊ�T�ޜ��5� `Am�����=�:��\g���eŰٗ��J���6�{�������ch�V�Ѝ�]�&z�/�~�-�]�Y|�u���g]	�>�$[k7���x(�O�I���[`.��QDu~��Х����|Sn��_�V.�y&�:����o�h0C�	I}������ʺ'F�����s��h[����or+����L�X�{�&k���g G4��:��B��\q��yg���m��`�N�A�j��M��ˌ��'uA ���-X9B+�O���A^�ۭep5DⁿX*�� ��>~��7,[��$+Ŗ�a���W�<]�Nt����
h�.�N৒8,��������SZ/��_�c3��N�|�m`aW���V��L3͊#>�ܾ��-��j#Q�;���Y��v�����:�T�hJ�~np M0Ɛ'px}���R'��O;�D3XL0P-�'�#gxR�k�Cu��M&,�f\�J~�:P=AWdN�\C����Z�G�l��N-1�`"�Cg����g\ ��B ��r�7~����Zp���᱁V֝��(�$�]x��v4���p�T���a�8W����/����y!h+��s�l�L�ޛ�Cti�y���4g�h^nuE~�$��>�/��du��&)¼VB��U�B� ���t:�̠A�E��iy�| �8��Pd�'8t��1���y {%�춓ݴš�n{�
^����1�6���6�+�O?*��HQ���8~��#�Ⱦֹ���}BRǡ�g�U����	Q(h<��Z�Ɨ�ن�آ���-��:��0�����up���I�p爆H	�cÚLx�f���4�G�UI-�͋�����O�xU�=����0h'���,P��e��>^��Q�����ʿԡ�v��,��<
�i~0O�Ґ�B��i>M	?��Z�+�׽L�Bc�����ho��^���,6��ׁ�(�Y�ԛVu��R����-Jk��{���U"e�b���+b_�yՊ��.i�^��+k����|��!- �[����p�M6��MT�}�7#4�d-@"�����V����eLY0ź�_Ȏ��s��(h���b�L)�-�����9B~���Bxߝ0�3�l�O�(�!��i#����%C�Z���x����k�U�D�&��M�7��k;�\����G6Z�����͹�u7���E��Ϻ���~��s�s��f����W��7�㍿�h+�x���^��Gb�?�C�s��e��s�@e)��i��xRo��DP�~g���2�����]�r�U�*`��'�|�$���&�V�Ӥ�H����!4"���5	:LՅ��N�qoihP�sK�ܠLۋE0��8���mĹ��]�a��Ix���޿|kPw��!u��Ǻ����Z�1'�pNǈ�M��>Ne��j/	9aXT���E-�)�Z��o�j*�ec�]cB�ٮ&PMHߓ�c.��%x:Hn�	���9�%#��<@�s���v\]5�����]'ey�ýP�wMb�̔H^�VIHJ�+�#E�s�k�e,&������,�l�0G--UQ����	�w�l���p�ݗ���r-��a�c:!��p�H�v�e��s�x�h2��g�+�xo�Yg�Qѯ�O}� ����
���1��4#�f���2+���+?߁N���#?��J{*����p�q~g��,�P�Uϛ��9#�~Yo�\�\�ˤ8.����.I��"��1�O�U��U��jZa-ǿX�
��>��nd&gfgLV+�1�W������ak�,�[����pFG$�A���8_��-7���P���T���j�Ǹ���m9ϥ��P؎�g<�<c�T����ݮ8Dtm��QfMW�w'�)��ã�������oM�҈C^[e�F(�ڴ]��v�^�Ø˗��{�>q���u�ܦZ�b">�عW)�������5;��������A���1��G]�提�XD|e39����W���'5�!T �n�'�7�����X���SzȼZ����MH-�z-��r�G\I���F�S���E.��"w��E�z�}-�w58��T�7T�X�[�f��*�9  |*�}f�2��, �	�H` au�i�p�����T����3��>>yx�$�p���I���^ߣ�����X�Uq-�$���`�-p�z4k�o�(Ϳ���g&��|��Ǐ�ƀo��2��7ط�
[Z����7{�Ů$�_YVT�.�[ԏy���o]]��t���ʨQ��ć?�)�3@x�I��'4J�gf�ׅ��\S{�%T��6�bo-�?	�6#w�z��1"�Y<����V�ko ��%g�ԭ��?��&�����㳸��u�݅�����9{}7�5�eh9:����d����G����ѵkO&!�p3��yE]��BǸHu9-r�V������0��%���	y8�T��9��שf/C��MS���E�p1�:$UypE~\:"���u5��d.�$^�|y�����K�	36�?G��:DXȯ��w���?�VHh:��t{����!�m{!�/���?�T9�_�Y���\[�k��뷇%�	�z�C2����1@}��ΊM��Hm�zf�=�6�H�WvA���Yb3��Gx��$��JVFG苸q����n�6�r(e�Ԃ_/񘸇ܲ����� g�5�����E
4���|*���u�E[2�"����Ӑ��D=�ȸ���lW�9�_�e�U�l�c"�#��g��/ܹ~�G��Z�����'=����
�eG���qb�D����%���&G�!��!����¸y1�(C��p�ˁu��߇<�!:m�6�
|��ك����l 2%��������׮b9���ִ4�;gD-�V*A��Fb��$(C2O��OC��&|}���*es�
m���M�]Yd�<�K%Ɂ�=2}J
D��D85A:_���qJ�M|��Qs��E���n�π�R?�4�ԗk;�anl���u�8��w*R��ܾO]�f��'�o)R�킉��Gd1���h�����d�ֲ�!��
ῲb���`��;���e�IT���ɼy��Y.�����^o�ɷ�~�O�:LB)O�F���K��(Ib.d�����>��3��ā���C��}aξnZ�,Ow_0� �L��:���J��]yƉُ��^^vm:�����Tz;���ҕ�j�A�/�eq���X���CQ�y�{�q�P����P��\
�k�i_��\v��l�u iPm`���ݻ�
}}�6>�]�U	Lp�P��OCd��M'��p���dtnO���D�}���Y�����X*��W����2�C����-����h~J��=�vX�S���U�쯱bG;*�:��9��,�ϰ���2���W3���H�P�Q���̒�O�{�Q
rRi`9�1�HFC��⩝i�kl�x�`zK��O]��*roFjq���|PrI��Nc�q��^ڦ��
���$�ܨ�.���dbekG��b�C��
���G����Ӣ��Xc+�ټ0��
�d�Zy����3霅�XjD����k�������S�K�8�X1�{Rw:��b��� v�r�p��2�g6j�`��Ҥ�u$��G4iM�.�A̘"��%YYYAa�K�XM��Q����B\��-�Rj>8H	��63]�����hX5�����_�D|x��a;�*���pU��p�ǪL.����J����������Y�2�y%���[?��X�7�}����J�-D�>����d�m4�h���
�fS�(���0H'�@��w����9��>�C��֡V�vͤ(��0>��UU,zL;%��ۆ	����I�N�i�H���Q08���5�o����z@�� �̚��L��0�6����		Ǎ�W `y>�~�D�@8[���ܤ1t�r� �=�&ޠF�w��y�o��r~Q�9c�QX9,�S�Ф�(45mp�=��"�&��2Fj���H�c���&ˢ�􆭐4�pj�<i#��/�4_x#)f�p�&�-Ó�i~�-��sGv�	^�%��uo�@O���@��3S{��H�0Erq.��Oƻ�F$+D#�MbP;c�)�]!E���HqݱV�	��_V�����Je�}i���T�Ț�ӓ=��z�����k1��q�Qr�����9C�����+4\��CY�C>r`7���t$ܸt�:�L�x�0 ��3�;Fe���b[ŀ����ҧ�[��j�j6�t�g �9�,�³�2���6����|j�}S��(����W�,Xۧz/Kv��>�sȍk��|w"�D�B�����z�WΒ5Q��2�Сu�Ĳ���$����Y3C�8��7��H����X�SA%�\�TQ���]����"I��`?d
��ع(I�yb*� n ��$���6"2Vb`d}Ue��L�@�ڀg{1MV�5��K5��`���/�ӰU�@L�&�jS��8��O�H�v�R��QCo��5!M�yBGA)8�`�?3$q��2���6S�p:��#x��Tؒ�ҽ���T���&ΜSm���� ��0�N�с^&�J���=	�Pڿ��`��kGۡD��Vd*����ߡY���]87l��D�*W���������5+#�0�*b�X��	�Ń
��<�0�L�D:
��?�bTtˍT�^��B�ۛ"Pm�T�ySq@���G�e0:�
�����#Mf�(�M-'WZ3��bg������;��w�r�^U]XL��EdY5fn��+r�Ak;�WWՊ�+��FuרoKb���bx��n%ݧE��;���N	�z�h�����+bV�?��X��O[���n�.5�%Ga=:�}���5� ��r��!��9����-[��
v�u揨���ex��,���]۬���u�[�G���e���k,l��/�V����76�fe,�jh���f]�=[88G����JI{�N�Ѽ���==���/ hB��E�G�!TC���(2#�54���ED�t�FI�<�$�=}hX��p��f�+�jn��Vf��x6E�-�{㱼��
͝M���<0A�0O�)�s�S���̶s������p-aX�#��M���"����_�퐆߮O�P��sQ��@/U�Zw�s�mE�m�U�|��0�R�Ra�AX	�("����[/�U��'�$%B?]�sΙGi΂��}�ϪNZgs-m�4�MLD��6�}%s������ �Mۍ�!��B���m2�����a�sk�/0[�.�^_|Za.��j�1�zH����b���;C�҅9y�.Q�"���D��N)�a�9�k���ᆥ�����]@��u�gM�H�Qt�	��V��~�F|9^K|]�$^��sn�`(��lY��'�q�ߠ�	���iؘ�Vl�R��9	P�C��J�������uz_�.z�a_��i僮��k7�������K'�m�(���8���U��ӊ� nw��Q�9h�Xr�"ܶ��z��O�L+u���%?��ύ�y���S+7��V �Py�=x���c|

qf˭���-�#o=2hX�טBȡI�Bs
�x�	�]ɀ������}���A
��ptu���Z� 	4�+Ŝ��L��G�2�QA�Ľai.N�~Λ<���_ƚvZ������-���f��3��n�����U8�ǜ�/�rq,�)fU=����r%�J���+�w�p䔛�gia����=^Ƿg��u�^��q5�Ԉ��	3k��C����	m힖GȡճT���=���y@-��J���^z��adϷ��l�+F I�!�G>%�s����5���{TS�P�W���U�ޝOܧ���[�����ׄg.��k�^yv~�.��S���A�����] GI�V�z%J��G;^�(v�^H<�B�k�#]��$N.���$��Φ�Y?S頋���I�($)~�w-t%T�&H/��47�?|�q=O:ٙR�|F�}��ɯ�9�C�/h8�P�[�i�8�=�=T�}pӕ��	�T�{���D�����"�6�2n)�Q d����p����p�rx��|ȼWg&uo��A��l'�њ���+���n���'�q���*�k ����U��DC�D�4��3�Wh��d
�6}�W�e�{�c��RHy6r��!���5U:�P8q;����f�R_`�hH*��)��(:Y���[�Lja����0v�+��ǂ�q� h&�R kq��
�Ht)k��
�J��"�3bݯhTҚIS��x��B�*7���[j�覭��U��J'#���v�=3|m�!_��w��A��:,D���k𜿈��rXC3s��nU
I�e�8����{bj�F'���z�R�
�oW���]�j̼��9���G���
p����{l�X$��l=r�Nz�����7��YYa;��۫�������D���������k{+��������3L˓WIŃlg���L�p�+� Zb�?�e�-0����m�)=�p��J�lD��)M��l�fA5�����g�m��ߑK��`*��<ß�Cݣ"���O��A+�����#4w�rs��u�K�� 3��t{'.i_@P0��r��R�#
Rh���nwÃ�F�����ߦ d�N�3���I��	�"G��!������c7���av� ��쇞w�%�`�b�,���^+�C�S(N�������b��b���"t5�}]��\��wE��4`(�u���'�e`D�
�=,<�&.<�hݲ�Gy����
_����"S}{��c#	�wi��(��ซy�Qc��W��4|��p8�j4������8_�m�Aҵ��c !�g�ՙ[<�����|�g��'�p��e@޻�9fo��	���Ubz���T������
[.���� �������r���T�N�%�q�.����^W�����n�~�b�G���sYJ���Z`^5����:�c���|�u���r��v_����ٵ��V9Wm���W2J9��&75pc����5!Ϝ'NQ��5�Z��;T��6x"v6�L]���(�Z{���3^"�r.��dȬY狳���[�9�Pry��T1�e���SAC���>��d�q��E!��?"f�3`i�����50h�s��"̴cJ��.�/ԯ|rƶ�9cbL�=t�-m!��Y5���~����h����=�Q�82x�cC�؉}m|A�I�"֚�+��̫#��0��`K�d�y��cR!�Rh1�'�ֵ���9c_24Be};�j/�5�!\����a�� )b�R��_���y��� ��d�{(��kj�t�f�qi����Զ�e�0F.]�k઻1#9����/���T�|���'Q&I5�l��p�|;����qQ}��Vz�/3W*#
<Ո��f8���OG���Rx�Vْ�kv�t}:�zz^Ղ�Ӊ�u����t�l���ߋu�xb �:<�M���v��ZR��-���M�4�;�::<�Lyc.�"GU�zr�		�(#�p����TEy1�;�Y�Bj��|��>5]m�hk���GvuO��M�3�=÷9���n�j�4��W�%�'ױd����x+���f_�����x&��m�f^qg��Q�'n���M^�N)����,��ԍژ\�j�$[�D��X�Ù����!��������\�RC�L��
+4t�P[�Z�$t���' �'�FA��]PV�R�C0a�=[ e�҅4����f���"J}&@��� �z'z��/�'�5G�!E`cH����?��@�be��Zc����k���N�7�v����@6P����n-��~�����T��F�{.���A���J��A�����>=�pY'�zY�%���~���k׾�`O-Ѷ���K�ގ��h�Ps�`Lʗ���=1dF.3��є����G3XZ@~U�R$lj�{62�� �b�j�U-;�~EI��n�I ������{���X�-�	}_:�R֚�ܮ3�m��j\�uh�l�0f*��S�����7�Ͻ�Q<��G����?����}�R�R�i�zZ"�
����+D��l��)�U��H8z�v���^,i&P.�����������k�X�|� ?+�1����t�U�>��!�G�﬿������o��x��lE��.�V)�/�^���風�{ �'OL���)-g/ڱ�+\�:�V^��R�v�3�o#���b�A��ikY��0����ٰ�^��8�ttd�<�a]Xٷc+wb�yvMb��i�������Tp:�n��3E׸bN׆�s���PD����U�K!�ƞi۲�c�Ei�[�F�t�m���fA{y"0�sB� � �Lm�Z��ue�����TS-%�����I!�D�*ݮ���'�U��U �]]t 
O��.���[#3\�g�1��ݗ��4G%fE��G/�;S{c0%?��=�!���9y�=7/�)-���u��p]�����Ɇ����A'FAq��M������l������?g2����h�w��a >_�S�1,77b�b2쐫�vЉ�G�l�&y�qv�%����iރ���!�Ģj~���E �5����g��o�g<���z��Ĵ����d�ԡ6�I��m8��Zʱ�^E�GK�9׬$U�HאQ`0m|��߻wLn)�BR`<�Ʌ�x9.��ꑼ�G�x�ags�c��h��z
.��53�d{3�0"Dsl�A\���T��W=��|�L�%1�ϧc�:kժ�!��󘥴 �/8��s���ۼQ5��������b�((�E��I|,����hw���F�Ȁj;6�PӴ���<��hZG�qnhX֑�ft�A�5��Ƶ�]�毱��>�Ѓ�M�Rw�}�1�c�p�3�6\��d�`Ȩ��
�b`R�?�5��Қ*r�r �L��ľ&#{�_&��sm�fz����h!\��*���o`���X��-I�ү��O��D��T���y%U��݂�]G�µ�O�q����J?w�cZ�[�j+?v�(��7�5E��{hH�Щ��+�s�ؼ�	d��&B�N:j]a����b��h��h���e��#�)giB)1K^_Ns�E�l8�C|bN��0�yEL�B?{�N��J��|m�P��s�@������9=Z V���F���r�gg�)��5�W�Z�hU׍��U�z���/��wh�5��-c������qh�O )G͙a=: ���@#v�̪�|*��핸��P��{[�`l�T�6��M��۱|1��f�����Ёu�l[ɥZā#��m�C��M����2�7y� 3\�+�lnoJ{*� aW�U�kB/��^���H����p�Sw­�z���?�/&3���\�_e$��j�g���*{�90��P��6�x:��M%1�����9s*��sJ��c&��= KH�ˆ��UX��4+5x�j�b�)�6n����c���K�<���]���uj�)H��mE��w�P�(c,V�{ԯ�����>VeI�߲͠(�	�`�.��a�zcEvE��P���R��L�͆6R�M(�)��u�-4XZoi�[^�p���b�&/!d�&K�^��,G/Y�Ի�Y��XGI!5Yxmo�o؏5Y4��]�����M��q7��5��
֢+� K!qW��F�Rٵ�+������KH����z���F=�\jn/Ȭy��D�/t��p/���Z#)D���s%�Y:I���n�a�0��YjEa�c�EȆ�L��!Y�uT��g�h�p�ꕺWtf�ܗ�z/˻�L"��޶K��V�Y� �-��>|�^��J�&b�|VR��n�*�y�U��j۱>8�5�%!v�����8�5����K�
�*ګ�<ؑ=�-�C��0>�×<��?��~B��p@���y��;љ����w`��&-ݱJ����3�lTEw�p�EEp���Z|��I�D"0���>}�g����Fg��Yhѩ�<����i�t����VG�_rR��L�~��
����̌Q�-[�<З�ׂrΤ`�^��~���'��D�Ê��
$>�׸�5Y,m"�]:MO@��mI<��u�bR�odr���~�Hs�u,�"�Z��W��| �g	|, 2����Hi��]�1����j��j8����A�U�Q�2n��B}	���~j�s]�������M��ۏ �%��b����6�U�s�b+�=C���p)�&�8��5�B���)d&J�is����A�H�vn�� ��$[͇{�ɋx[�]k�G�4�x�1 �G;��cf�v�H�aV5�"��E�%��.�,����g@�wĜN��Sϔ�ji[��:[� � R��g��'���H�G�s��~-�o�ӃIpp]�l�жO���m�����a=�����=Q�d���*݊����|G_+�E��F+Ղ�/��� 
,�B��L<���&��f��j�Y	��qj���G��BF��rv!�y�7�n���ǥܲ�1A=����,�|�U$Ӌ�V@(��B�{���"�!�y?g>��Ҕ���<Z'�f�:媷��A|�o;1c��Wց�B�q�J�.��3��?We7��m����w���j�����ο�PJ��/g��8��U��d��
�ŕF�z��Z�rf)0��J^9�M��O��I��)����A�j�4/;%����a����Y�����@�%�O��;�iŰ�JRx0O�B?g�qNJ�6���}Й��ԹQ7D�%ﾖ�ݶߛV8�}�:�j��3� �W�c�r�h��-���1�?�g�f��i�Zw�`^�����ݑ0�8�C���$����?@H������{)C��wj�p�ۛ��U����Ga��c�A/�%h Ytz@"�Bo����v�ct�OH��q(Wû
x4~�<nUF���R��̇>��8�E1:�w�f?e���}n���a!G��}�A�!3��H�$��ST+���G=@����DV��|)���}��3���I�Q�ZΑB��+�K�m�I�I���-"�k�y�k��$h�6��8V�B��]G����Ji�?���T��id�⋹Q�$U��7��`���?�g�\�K�/�.��7��|Z�� Uū���1Yl���1� ��]O �#��{�{�!$0�ZY��OѰ�Y���{O��Cs��	�wq��zYs��T�㤠�H�D6x�6�!�ѫ�<��~��_�Y[G��>�dӵ��/f.aG2����c���[��-/�$#H;3������0��m�g��Zu��������w[1e/��K�����E=D��F���w!g�*�G-l~f���S����{����s[���o�h׊���B��c�;�a��`}�+|F���g6���p���GLJ�*�q����G��7搃�ٮ����*[y"���f�q�]aU����-�B�{y��u	�,�n匎������KC�3��XhZ�j�3�R����'7�{����W	�֖��`����J	��!���YZ\)^�:���z�������y_u�e��L��΍0y�T!́������:[k�mI�虣J��]���Ҟ��We�j������y#���Τ%sS��'O���
<xl�h2�_����b�>2٨�����8	B�G��w�SyÏH1��GU^'����V�q(������'>��_��mm����]�]@,�40�*t���0v�٤�)�;�%�Ϥ_��q���qspvRk��8"bC���8礉�DH3{�U<��P�C�|��@w��Z�R� 1W8i�׻���9U��GF�����mx�-������;w����W��X1w�h��1r�Pf�f�>�c��_'��/�`���MT[868�'�Yҽ��QCf�����1�	��݊]�B׃XKu�
e۷Ywٴ#�����e�|3���ȥ�e"]�6����T�}�!o��
Y�e8Ο	�ޓ���h���*��%�37����m��o��p�L&��E���ˣ�ֆs�`qՅ��̨	R
z�qa!kz���jܩ���[?YI5Z�u\( ���V�&kkeT�Q��+�g��8Z�#4�0jxs���^\؊2���7�����\b@�͂�N��L>z�,���)�[� 5{R��k�������j�kN1�I���~��	|' q���(c��?�@�MN�YKP8��K�5}C:�\��-*#����+�$%G��g�U��;^��E������:��=)����/��`�;Ni3�C����g���� J5�(���J�ڶ_�Ɇ]�c��y��Uq�*�G��2g#��g����70�4bO܃r��{`[\���|	��E��">�F*��9�~��E�d��Zϓ�)��93�E�wo�3�����3Z�9-����,��p%0l�11g�� !(b�]�O믲�@#�Ix�;�\�)_�L���$,/װ��1��( -����sN#۴�n�>����!(�3'�H���)I�"�m"8���o��(��_J�u��o)$Wc(�]����3O��ʓ�]Y�vg'L"GF�N�8x��r�³JX��/"���>� �1l��Ƨ�jU�"-�����n�R=&)�OvZJ]�O���|����\�*�hWuY���> +rw˧��v�~���l�����M{��\0�T��W��	�C���F���Wɺ�R�G�w�^HC�oT�A��*m@�1�6O��ˁ��<P��P�D-;z�?1VpHĢ�]Ҵ���s3"19ч�
�#��_���S<卑��v�j��YaСS�������zk�BɕL-i_ �uJ�����q�\O3��	N�z��C�$��^��d9É;�Ѡ�N���65��B�i�rP��y�8XnZ5����2s5uW彆��X�h1�A?4W,!t��P\�<��#T�`b.$���׼����QMtkn!N���4�IwD�G'�b�\�9��	9$��cIp!��2���W�a10B�7W�j�4y��@FQ9��& Ρ���+c|�5Gst�0M>�g�񁨎������YbS��<'��N���V�����s�.�#�:*�	2�]�д*�h������U�L:p��}��Ic��;�K�1��?�/��԰����Ң�y�,y��x�{-�vb���P�5�^��%/} s ��M.�*�O��(�@��Hئ,���O��Q�"j��~�,i��k���1(�=aĂ��`���iq6��s��Z�Y�aQ5�ָ.�"#_�
�a���	��Jդ2ʂ��z�u��*Rl�O�_
<��<1Nb��Ca�g挌�⩞G�1E�I��P*:�`G9ti<���`зg�s#$Y�8���S���R�(����اc��:��ﰨ"��*�&h�"+��\8{v}hr�]�NPTd���aKۗ��#�O�E�Ճ�q�� �N��7�߫}���i.Sz|�YU�X"�坤GhR�/浹��k�ʧ�=��I��p�
���k��(� �!]���ׁ�Эz�D��@��� 
�����W��g�=�-;��R��;8���*��k��R�75
�@��O����k���)Cikf,�:���PY�t���f��7�}�'c��t�N|��b�a�����Hб}��O��S:`Gt���\U�]m���1^E �L���P�HA�&�`|�L�D��V-�Gѭ���ƯS�������^ -'��m�O�~|�������y�����T�S2iRD�&6��p�t���󌝠���B�JT!���C+kLC�;q$��&c!~��;z�Q�/�fi\<Z���ò� ��	�C��e>����8�Z �%�v�5�����T��p�z�%��� ���)����4�����鬤��1��b�Q�R�{P����	4�����\�Tke������o�Ņ�������;��EH�KM�|)a�Q���3;f�������8���i]w�Q��� �W�8ʚ�9:˼�Nb,ef�o����5�P��������_zF`F��[m�ֵ�YK�'E\u�>�zx�z�J����~8�1/��U]H�6V�����5"|~�M +�qo�J���߆"�rک#stȀ���zB��>&���_o�cYt���-�U���1��B�fe+��F�����bYY�\@yD
�]_9{�?��s�P�c_�WA�:�a|�D�m(�X����m9����h�U������O��5�b��j��Ȱ=��j`V��x_��y8��k�a�*o�v|l]�
�D���v��L��:P ��ܫ��.L��K�G������{�gD��[~tO��k�2ֆ2�sn[�t�>��\e�0��Z����Es�q�
v)bU��w����.���F�����M2� �G��K,Um�Ü�S{�P�F�>;�\����Fbf弣�+�@Ȑ�""�Q��7��d�};�̝�>^_�Rz�a���1`�����8��ƴ�2���pCvqB] ��"x2\��ѳn�!?TM]S�7�#@��S� ��cE�Q���pEQWq�٫��j.��r��w[���;b���R�)ɢ��q*��ƔTd��ܣ��cf��}�sԍ�p�Ǩ��W܁hޖ̩
�xh�P��؁ s	�vf׬��l�8�0�j�'.��p��+�ٲ(d��(et��F��~9�J��ɒ͢a��6�d��L���I2Ь��FfGzl�}+��p�yum$����tȫ>2*�t�%�1�;Q�9�,�l��a������o�̞@0\?�v�����H~�7xpM3~Y�tm�֡����������һ��)tNד9Ib�!���A�Iu`I�µ�@0x��|����#k�߲�5lg0��	D�6I��@V��h��pl+����� PsS�@R&#��]on���迴�A�M�T��l5y�ϵ�\�j�hw�ۺ���[q��
���@OW ����L�wE �eفd21�W:"t����L�H��IԠ�! ��f���!�W�m��^Y��
U�B7���K�Ci�!W�o�/�ЦA���_���"�/j�qr�~5\�66R��͆�=��o� �z����G������[�Kc���X��Q���߂Y��~� @5H'qG�:��U��E����E�����I-��9��$,��1Q�$aV̋=w��w&�߸8a��S��������F(H���%�p�0�>{��zkA���pYg�a��T�R 7�惰�Y�GD�?b� ђ~�� 2N��REK��Č�e���[�G^�|xO1[�?�c̳�rI��I�k9�ƒ����g$�H�8��`Y쵡ş���}�	��C ��Dr��ٲ쬀�c.bZ��)7ηꑂ'�{up�>��f|Ec���Dp	�.����|�0a`y��X)
󙩻�M�9O�޻W�W�@us�_��P�`�J\�4J+���f|*{�Eզ븦Mf��U]g�MFXI����ݣ��f��a�d�t��Pz��j��A�G��]�\yI�_`�����Q��ц~:dlꆓD�4)��^�O��Z�]@�ho�Yb6ދ��ݐ,��7���|�Rd����"�X���a$��d�t��#I�%H�_AM�%��h0�6_:���R�u]�FB�ڨ�l�A��0���y�`$��"s��	./��b3KW$՚j	@x��Q��<���TL�X��֙x�z��w�R�A��b����'M��^hN�Գ^��u���$]Հ�]���[��N{�k�67��b��c��B���8-pӽ�K[�ul{��<��C@C�],�6�
�MJ����\pq�&�D��:�0��b?�;W#ڴ�<�u:p�\|�|��h�C�e�m��cyO?ia��Վ��J�$`��tś᤟C5��of�E��xki�-A]�j���gay|�E遱�/$�;M�]{�9��8�%�2�m�Ҥ&]��~�69{�&���E�=������_�Rx,��N�4= I��v �[��EZ��hvoDk�@Y�!��-����{�~dM���"D�Ș�%"ɐ��CY&R���0LR�L|$O-�L��NF��B����l�RX^�wZ+��l�'���,��1��`Oj�ٗ!_AI���Ġ�	.�d�t������ ���V�ݷms��<5tKT��0�eN���*��-J+e���\�L�(�0Y�N�G���n!6]��B��D��K/Fl�d�|�u��:��:��*��:��R��|k X�͞���:O01���+���d�<�Kn��%ۙ�ۑ�Y�a�&8z*�_f���������.�b��{��8H��kF��"�?-��shBk��a��&���Yi�C��U奵'�9%�j�J�{�
��R&ĥ��������#f��-z������y���(فz�D�G�MI��H�*�ģi�E�+_Ah:�#���:�i.�A��Ȧ�m����T�
��Zq����%��J��V84�cm2C�s����e�Gpx�I-b)Q����x���ηX��E�!�o�X�U�t�^��81�*��,��H�<�͝"��ɌU+��`���|��\�JD�����j�iz��M];�hQ4J,�����B���}���#AGZ���K�GEw^�>��5��J�[	 \��N<����B�����A���':����K���ؤ�2�_��U��xQ�@T���*�����&�PD8��R�(f�]@�op��(��e>���+�ɱ�5.����؞豳�����ڣϣ"����Sޢ���C���:F�|�_{�V��P6���L��i"����*ԯ�˦e����I��r� ��N�ͨi��������8�E[ؗ��e�F(�ɀ�vW��ʋ�����a\�w`鲫�L���G�z��+�G�L�����i=�;(�H���{�<��W^�c���p������3Y0�*���}ךN��-h|Q�����@k���h��"����o	#��<qN�h�g%,�Ϳh���3��>?�qkSB�K��?���X�����m6<�����`����#ʡmqWiZ?@��M�H>`%�ص��8f���� ���Y8_��1HD�w�E����jd�@[�ݲܡ�`�!�6Q�4<O$]����S��h��II�� �2�"��y\u��νmĵ���h�R{m?Zn�L���+�	|U�"ײ�\f#q��s^��
�.�L)�Eۄ{y�Z�9Ô3[�[^�˘�|\�#�8����?��^x���k[G&��
�U�Y>�Ln�Y�N�nN���w��ԡ��I���źCY�L���T`��T��bh-���Sm�������ƨ��6g=n� Z�GC�� #6��Y�n�A���
p��t�ba�7![�A��6���{���2�"/'(�?�<4+���<N�Gm�j4m>�x-b"2� �@��b�Ӛ���{��c鍊��Gq*S!�-���
X�B�i�/O>;Z��U��yo4�]�є����iII���Br��tX��j;��r��\0\9]�/A^��#P���e�Y�2�B���G�-��k�\��H�T''�$�lx֔�����&
�o�0��b���\�
��D[�Hs7�����;k�s����h��z������E�V$ȗ�d2ɥ�N�8�i �����ѝFx�Ά�l"�7X��Q�r���S��?�Y�D��!
C�/������sB/��nWHv��
�*4ꖰv3��8gu�{P����J���O�	��.�'oh�DHˋ�z5~1]��,�EF_:�IE���c�4"��KܾI���f��7�.�|�DmHGi�]�C�U\"���e�~tu6B�B�����w�ӫ�I�u
b,�h�e�<��
�OΒw�?��S�&)�6KM����E`8D>z7�V2�Bn���^��vL���aڱU&̶������C���u�;㬔R�&�Gte�[�Ow$,���Y���4ݤ6������ ��ò�d�"<�KԠ����)9��0��ڮϛW�#B/��hR-���b1����x\�]�g$�D� ����\����`�6�/ƇH��4�LVjQB����뎠�Q��i�TاͶy?�ǘ[ 
LLqG���V�a��Qj��J��0+Ԯ�>p��n��^�Ei� ��!`���C��"���0R��-P�E�]�'�?D��d��L`�0@�f= �ɂ $n��Y�[�R���A=�Kb(��v����ٌ���z�Jv%4�����G-S�Ѳ$���c�z���ds:� ��������H�M�X��ق�K���"~�X"`'��d�����Zgkxz-01jCEs,�G*�T��LxN��+*'2<f�N��ޣ3��y�#��}!�O�X���[�&?��xp���it���

W?N�J3C�'���u��]���Z�+=�[4<_AFZ��Zkk �$����d�������B�h�§���t������|w�8��ݟ�U�/CG����Ϧ�ԍ_K9���,k~K{S#]��Sȥ�{]܁�d`Wa{����֢ߴ6�e�&Q��_m��t,�Z�1D�Iy>`�@�H�ɤr�!n_[Ua��(�3�/���bk>M��U�$3W�٫����K�N�L����/�1��X�na�țg���`�Ft �T���KLⅷo����A+��l,��lc��W6���+1���mL�;q)ds��y+wEb@A��d�8�;���ylg1ʳ��t����?�K�~o�Y���M��r���Qzf腪�H���X�!܋�X��OJ*K!���e��0`f58�%�����E�]Հ�1��]�����՜��Bz�3-�o��uB�Y#RxT���4ؼp>Z�mz�Їdlv�ҤT�Gt�eԈW/0*|�G'F61���->k`��><������Tr��8��fN~ ��@Ȑ!��:�~��_K�N����`k�����-q���z�~�s�:'혆<l����zU R�=~�����*���cD�Ɲ�HNˋ�g����;�bs�s1x�K�Jͬl�ږ���z���}�̡£�>��O܁�E��5���x
��ƹ� d;!�\x*EՊY��>�ّ���qI7�
��>dJi$wd��/q�*�x<sM'�!H���@�I�(>�
� x�d�Fm�^t��������`D5���ȋf��0:�vY9Y��]��bbؤ����q�Y��Ӏ��ӓ��RY3/L�P�~=�~8��'�vJ���v���]�+3,<��%2�l���p;d��+���m�������Zx+���,���س�eF�ony�$���1��P=lA�}լy�z2cHJT���&��$��Zyg�X�]�},�Ë%�ӻa����Hg�U�X��;�^<и� ��9�R^r7�*I�|NS�kM<OIQbkS�����\Aul�Im�,\�1���c�H~��A]�Y���y����V]���s���J�33�M�l�&��z��Z\��B��^˾�
@��Dru��Ki5L���l%v)�N�����'�rG��PR�����jbo�̇���,�q�w7b=<�_���AszVK��4�/��n��J��'�4��t�d�e$�Ӓ�~�v�4�?�L%%�1+��) �$ke�$�������2!�?��QQ��NW�b��b����~%*{���x���2�����Ǟڇ�*\w��#��%�"�3���y�J"1|y5�����Z�����L�+��g���nxͭ�ܽ��Y�.�[Y�6��+<���<�X���ڟ`��R�4�d`�c�x�e� �0��H`YT�H�W�2�mۍ��(Z����o�i@d���z�^�1�U���B�`�L������>���x��zh�3 ��[�sT���ݩ����׌�K<����OP��t�>mT1�1[c�cϟ�
M�� ���k��OԜ�opoLm�z�h���"�M�=r���nA>�E���M�>/��Y��J�֧1=/(��5�i��!Wu��Iwߙ��i����� gxb�w	n����bgD���*�����L�'N�m��;�ϕ���v�6��OS�*������BԄj�밥�ԏ��	j��nWE=+O�5���N�J��R�qj�컆.ghu _�q	Cx'#���x�Z�QdA��ގ~�bW{nϔ1�MC�κ���J��jm-Ys�?g�8b�
	��v�|��,��ܝ�l$S���	����g� U��2���+���N�dsQw�\�LѬT�g�WU�.%�o�P�lw���8*�OqP-g�~<�8R�\a�8y��1h����'�r����.���t��[Ic�6��\-��Nzy�mEoṜ/b�U#�����*��o�Q��Mj���
��O_�����<�9��X4;W9��S{�n͒���49��O?8�7�	J$^�.)O�?8�5a����Q�7�@�-O��A��&��� �LI�';���O.^�=���./f�h71��w������8&6�$���!�w>��D�|�jgѩἂy#jp�Z;,N�o�v.2��;��3�9��5�%
|sP*���ç��X_��ߡ�r$¤��+���
㩫Ϣ�r�;K�v��,���7���|�7��� �'B�k��U��5�1�էkq����H]�.�s	c��: ��Da��rI�^�ex� z�TۄPF�["X��!E�N��"5�ݑE?��}s~ڎ���\ّ���l�P�G<0�'�1 pU�DۇnO��x����Գr��Ef��κ�����`l~x۪��͑�Yp-��!}�e���醈�0��}Kq��~0*�2H�[Fѯo'[���v�`��$4�aM�e��_�����R�^B��y/y�p���o�։61ȉx���8��3
��ʘ2���/_�-�ume���!�{J`!�{�A�r�8
��t�H�u?�iL7�Ʒ��j�aB#RԲ����?H�(�鉵k�g�ux~�u���c�"D�J���#���:�@�S$}��������N��1���ǈCg-#{�� B�����	@�4�/�|$՚�c��x���&�y�V�[�9To��0��ѿ��!�1 nM�p�?7K�^a�v|#Iw�vG�{����@�~��T���#F.]�^di�n'��"]y"�f�1C�
	=�^tRs��]�#���H�簳���@/��%�G�;�,��m�#�U��"N�o*����\L4@�rG����-o�i~���e�ž����F�L/��'_M�zU=$��ۦF�O@o����Bp����z�,kV(�(��� �󬃇��eV�$�(�'h�y�0 �r�l��R|�i�B����m��?Ӛ�bЍ&���Fx�ȼQ�dۓ�
�G��g̈́�|z}����8RxX���M�y�paT�{�*����y�[����UR�<�!��#���t�T���Đ���zdj�
��E3歳Ҫ����,���6��V�FS�uvz���&QE8wD`/h�f��a\�>Y��BK̬G�>/��z��5RG
5�Ʃ{�>l���;���`):7��:Zҳ���{䰲K*5Y��b�Jt�z�������O\4�}��Nl��\�xG������ۢ˼�?�l��o�Vm��u��~n�2{"P�?�8l"�"��J� ґ�_�����pQB���f��QB�i�'����&�V�R�}|��cu*6g�῞!�Q_8�|�,P�1x�����y���e�aQh
�r�n��0t~��a+A�i?�!hJ�&�
����-ex��A�+d��V*0����[��=��5v�é�+le��ѱ�_.�� �.�`�{l)#��;����>o�.��~�0���P�t����j�@��ik��ϳ͛��D��7ɵ�P�{��=�`X�A��gd�&ō,���ZEJi�4 W�0�r���n&�](�m^R���ve�CW�YiC�k���OO�-��D���s�,��eT�d��8���(iL`SI�/�/vAm�ʆ3NQ�2�����?w��e��ʝ��0Q�0��NSl����Xbk��B�D�e�#���1�w�{��c
��$���x��$���Q|��Qg~-$#�΁Xۿa�)ͦ��<y�0�H����-���F��w���c%X1;�h�>!u���N�׊���K�,
�H&㛤�%��>k͞%�]5��k"�}V�c�9� e��%2<���C	���)��*��w��e����|-vH4ͭX�I��Qv�,��FL��:�tw�L���^܌��Z�q��S=�d�%���u��[W�Q�֊��+��Ƥ�L�D��N��³
p��w�íŦ.z��	q��82����P0�P�9n�����: ��T-�{�wC�L�>y\���Vԋ����-4.�ڝ{�]2kשnC��p�K_m�ALK��Ϥ����jEB�z���xYg'�1p+^�((>��ǌ�(�Kl@���/��qޘ��̙U��v�Q?��項%y��H2�����L>���Es�o�2�d1�����cHn� ���J�j��VV�B.�d3�5&�RZʸw�]TT;�-��bN�G͟Fx���hzȣ�u$4���4��%@�w5��>�bkK����ł8�E��3��p+����q!�R˅XqA��Bei<���Vߥ�f��;	����_�~W� ��G_3e�%����dh�p���Uy�IQ,��l�U��ehH��}y�)x�S��Hp;������яt�lj����B׌���"j���!ew��*��=���'�Ψ�p�ݞaL��,��U�E�y�(R��L�����3��X�K����4���#��rq�{3V�b��yY���a_�)7��ee�إ�yn�L���&�}�z��f ��r��5vr.�:� rrA�G�������!�噹ڈB��G�\��|>�H�y��!*���(���!�/Dc ��ߠ]ɲ��s��A�?e*#���E�ݿ6����WIk����m�h����1XP4��M�x����B�f
�<�����22�������m�i?�h�LC���ݳ��U�荽�\�|�&�_H�)ڕfE=��-)� ֥6�U��H/WN�j�O��@ƺ�{��WN���κ�����j�X��L�����d5��"&ճ(�l}P@	kP�ʬ�� �\%�ad[���+�	L���MP��9ǈ���IHM�q���J{��ΚR�2�m�@S<�΅��J�i����V hv!)���tw��W483O� W%�NC�I/�#�d�<���ԡAK�k���@g  �I����n��`e�դ?�p�����Z�B[��
6�&���|~@�r����=ϳz1B[���
�̦u��v�M<�v���(©��!�s����w<<=u�l�l7���S0A
_��h������[��\,j��/�i�Ⱦe�q9��^{��؈cЊQ�	�S�����~�)+�2��R�
R�,�SG,����&瘮׎� 0�>�߂&�Y7kAaN��ڝ�`߭���٣D�D�
�XtWrnk�A�c�4�NU����4a��*�v1���X��\\��n�H�e|`H:��8@���W�E���}�U��k*.7a��u���7<n�Ms~�2򭫊��[-��iwH�#�L�M�(��?�7R�l{�QA��z������L� �[l^�Z3!&�8�Q)�տ���"�`KlCU���p�:�L;���`���\��f���_=��}@��bl=+�������ʴ��&�qQ���ǘ���eŶM%]ȝ�*S$��i����	x��mg�
F�� ����R��D����mv����Ї��t9���K�,b, (�劙���N(��h&Z���&�����̈́�V;RV�� b��6!���6	o���hL6�ZRDm��qy���E�l5�P1p��؉-҈�TBO�x�Cߟ� [�ȞX��|Dè�����]��h]%J�0��O�ґH�FME�>	��[�͟�~��	e6͚�.*,~�M��^C�eT���w�n0 C��4�4��p4��>�[����8����\����$XWD"��
�D1Dؘ�3<s�)�>Os��kPNk�1۾f�ܥT2�ϖ�?$��%K��S��͉��z�rQi���HN�r;3�Ԑ$|]o�\��G��ޫ)y�:��泿�]mŉ��'N�t�u�����Z/��Fb(�V�v2Q̼{Y���تHֿ��9��?Z�Ψ�݃��OWn�M�k:΢��6.�i�u��F\kG���	��j��~���Y�{T�"��@�|S6�&ƫ!q�G�JQLݺ�ۍ�Xb��S�G��=��-�.;[u(x�����⪉�Ǣ�*�6]M^�z��T�;.�� Y��H^��G����ɴFkg����+�q�O��\����ރ�ï�S��#�Eٝ3)��{DlϼK4���t���@0$����S�!��ΛP��+� !4����H]�ź��cĐ�^p�悷���$ݓ]�|���,����[�ջw���q�~L�V�O��x�M�E���y\��'���k.:�9�8Q�5��tM�nG{�.#a��!�}�@�@KQ;4������&�,3c����[b��"]�J׍B�֧Q/���Ǻ��SQU�bR�fٗ�+Ġ�1��ta�(J���!�]L5�b8�=SZA`��^�k�7rS�x'�:�MQ$�[i��"{9^�U��t>?k�mӳn:1�rd	פ�"��w�4�a�N{��z�B[pL���*FS /���(�a/�xew�6��Υ�(ҝ����y�\��_����2K�.A�I�v.6���s���SD����4á��b>�G����N88P&��	�q|�=1�qe�*���ڌI�V�$�`cj*4��1�N{���P8"�B_��=������D���HQ@�	��T��V�;�w�/��f�<C"9l�i�M��|����ã\*��T��y�I�Z���C$��W$�7%pΨ���ip���NI�v0�3�ʸ�[�
���KA���&\nޱr�����)�l7��L�H�&����)�}��r� .��h~k��gKg��E9�ds�H�Bv��c�4�Y�G-�\`�o�C��xe�.Ҭ�#%�?��L��ß8A�wI5Y��[�A��
����},Xk��jg&I��)�����o�@6��3ãgk+�x�)�y&aK� ��P��Q���`����u�&b��*� ��<5�2
zT޾Q�����j&P�aC��4��ײ��ɷW����0��ɁZ��'6�������s�L���]���Z��Av�8u.����gM$` E��ݑ�c��	!*�I*��;�-�Ӽ�l�6dy�xP��q]t�V�%W�A����g0E��~�]�v%H��ҋmp܄�<)��b�:	��O�X�AU%A��|fZ]�h�M;<W��[z�+�c��γ�Ϩ�Ч��BX.�#�e�7O�= o@|�È�VZ�)ҁ@L!_ԂԵ�D���M���9t��}�E|2��x�^�� �?{:�q�� ��x�c�V��,�Kd)-h{��D���ON�Cz�ͫ�fҟ���ڣ -ش��, �;w��3���f�27��~JJP��n�g|��P��C�����l��~W��3@E���}�H����x:�1T�v�"�{�u<��
�-W��"�v2�I��U>����- �fU�����*�eP�0��m�)�w��B@���@�~��L��`|�S*�+v�n��[�ܤ
���Ul�t�|��8p�X��;��Nm٪f�``��M:'��o�Y�s�q���J$F5(��^!61�m�ׅiq�,k���ޓ|v:���m+Ma�1��m��/
bq��V��(���D�^�=�����]����	iʧ�sց��,2�����P�{S��ʞ)��b-p����ZH���,� �fF�������(��D�©CJ7�{in<�C��H({YbA��-��n�|�( ZT
�a8
2Σ��AK �k�ɒ3ݷ�!X@�׋�	T��ew��qT]h靵&k�|�-+��μ���|cQ��;?�(�gj�]c�5�RZ}��5�-�G�Rv��o(�O`�A��K���,䒫�q(�ۤ"�G�J�n�{T�&u� �ȟ栎 �K"E��z�O��m�������0�g�����E��R�t���q! �z�`����I<����#��xe^�v^8���t�\!O��v(�,˪a���:����6�	7��~[�$ѝ���_7U��J�*��q5Y�s�Ǫ
=
��L5pf����g�P�6�x��,��/�Q��:�ZAhj���0BzA����Ib�����d5^�%�E�О�m�YOp%��������І/�:��p��S<��IG:�4/S;ا�����'L�q����\�C����z�;����O|�~X�E��%ɖ��%IE�j��ڞ�)������$_�G_p5�\������u���<z��<!ï���{�\C@�1]�bCQǯ�-���w`�@&}��Z�s��]�l�&f��h����;>[Ӣ�r�k�3b,�t����\Rk'0�	��j�v��ņԥ��:�d�ꡎs��؂��H�4W~n���6��Zx7�Q�i�9�?�*�^�
��fvW�A�m�ܦ�#����'獵IwP�W&��a�d��[����TE��
�A�PF�L�>Ұ�]�i��!
�����:�m�Zo�����n;��0�%��U�ur8O� ���x��������֕�*�7��7�W!�a���?��X�(��:`: ��cܶO�E��VO<� �§���;5~x�_��4wv��?_n�sy��:l>��X�������-V/��Ң\3�ԋuy�@5�����'L�]4|�(��Q��Ŵ�{�8���҃7�;��Ge�EaU�]�V9�w���#G�hr8�ew(F�U*�;�k�9���F��`(��7ʽoi��R�QKC��!�(
�G.�0�9g��ow����#fO��Jq.>����M� �(�^R�Sm�;E���L���3E���mɓ�1TO�u�
��Z?oLn%Zg�Oc�@����j���*
E��~K�!�M0�L��i=�q�"VÅ]V��%Enk�kY��>³��GC��� V�*�|��b��MPW��VY�$-���_�G�k��� \�#�\<H�$��q��[q�hīJ���F�x�v�ͺ�e�V#��@�8fю�Tk�&�s�Z4!�t�6��l��Zx��ZRI�$ȅC���d�ͽ8R�ƞGk�8�=���=�{�dah�t!����7��(�>P���fd�y�N�ś_��]٪������k�$��,�#8��F��%T�@|��׳���׿���UT�,q�`��;CcW��SGL�t�W�k'\��S,���Q,�Sz����h�t�}bB�W����𥇏�p�<e0���P�io&9����R����u�g���(:m{���ȿj�;UY�Ie�Ĭ���[�����R�k�tR�p':M�3X<�I���"<fv	�v:�-t{&�~oo'J넔��
_�'3�|�� �o��J��k$"A0����!��*�*�ͽ�����op�|F!o�4��G�>�������+���P�����Pb�|6J����B ��Z�y�����թ�J��w��Z�b�E�4�	����F$��c�_Z��ﲄp�l�F�i1l��ݸ�`�>�l���<A�}�L�w]��@7�O�8w6?1⹮)1^�㬱L�[$N����7:��X����mG;��	f�_���$�����5��oQ�=�Vm�x�}� �n�&� =��Ӵ�Q!ٖ�V��6[�BjǠ�rZ#/{�������L�@�_ŷs�G>��O`�bqn��_��O�����&������,�,vX�EMє�L��h���g�c�|�ޓO��R~��&�d)3E�H&��O�NGJ� ^����v?��t͆l5������:��t���ec��K!���C�
��˹ ���ŭd��+�����ko��^�+��dc�a�?nD$����$���0�<h���C�5<�F��ρ3o��d��UEtP��m��j�hCw��g���y�5 ��m��r�f��n��g~iD����{�Qb{��ɞ���Y�h�p�����6qz���1�8�-T�r#�^�C�Ůu?�*�P�E�n{�����ybO@ɽm�l��j���i7�7��ƜϪL���X�?>�im/K��J��j��+�j68�(Q�1h��Y�-V�S�a"3/X��Nay��I�5}�@�s ��&8���s�1
�)���oT����G(�!���B���y�}B�@���E�Q�	�)���neq8��끀���kHk�<0��n)7�U������
�8�Ѩ�V#)`��	_s��%�^A��J����0$/x>���T�u0GpL��͖�:3����J�s�J#:�&�Ry�0�C�opUq͵$��%9)U$�Y|vY�E��]
l�@�?N���ʭ��e�(�����/�;==�S���3-�f�]���eJ��T�] C�Jn�r�cD�*�ԤiC����JP� N�L\��]���&���*��mVz��gۮ*�G�I~�M/����#�&��o{�m�y�;8 =�W!� [
X���<�EX�K\ԥ	�գ��"qS�,�P�n����Qx^��zU�}_�Ļ��m�Q@G����S�͛�q�Go{�a5U��:���gh24ளa��;�O�(�?�֕�����Hx�Pdatoy�*S��w�S0nh�� �0�Y�tK���<���vv� n��1��י��%wn��n[[}yņR�	���I�Xm�(i#�4�������.`)[�2�F9q�3R����7J�\��x��"1���P�e�J���������u�{��t�;���WiӤ�j%�����}� yMM�+͸��_�1�m�~՜*�h�2��ޕ|Ү^�ن��d�}���e��8�J�����)��}�L�~|����i9m%�B�^ȧȴ]s3�x�k�&!�R��	-��3�Y
%ɃP������V�R���)},>NC���D{n�ɵ���	�	;3W���zW:ojj�Dܿ)~!N�8�\E��N�u��3@�Vׅ�pp�w�$!IB�Vc�z~фj�U�e�@����C;(~�^Ժԇcs�W����H=��Pf�·��C-ٹ�CId��vE��J~����\�B����aS<J��N_��)�� $�1���k~�jKx._lX����|���ٽ�N8�k�t�㵓��v�	��^ȿe�d���n��aK)ڟp�niK8��g{6�� �q7LfY�M^ow�8<��f����0�d��Y0�U��s���sqp�i�U<�#�]�"3�g3�RzY�OxG-b����_�Ri2Ս�/�	X���H���x����k�=��!@(r�q��2��q����y��p�q����H�	ٿ����=y�yUJT���ƞ�%ʫ�t��X��9լ��Q�$����"�2 F�)]����w��ņ[������ZuUĎ1��?N�B�S�(�S�IK�և�r(�|�2_]�h>^	�{)S^�<����u,�W���LݦSQa@�3��
���G�˵����x�_E=�Ƭ�YwR�>`�z��@D�M��b���WL���1������ɫ[���e� �4�+���eτ���W"��Ua؃��)-��&��ޔb��ꗧ�Q�V�bv=pB�K鱊{T���2��w��������8��\��9@���f�m4o$�/~s�F���,)�H�`+h� ��3�%ϒ�y#��c1����:ʆjम�;ED�㊧�d$�W�%@7��3RX��������J�ϕnh���N��?�%�&,�=���MϥH�r8��OE&}���E\_��_U�z^
�6[����*?Zrf�1ە���� ?�����yEk&��B�0g��v�
�N�OM��,��V��d��*�+�IwA��k9}B�2fց��T�ě��NlZ�)#x�{!�"CN$2�M�5���_��>{�xS����2.!/��s�k�jJe[���Q��:s�/Z
<���^u/p,f�h��5�q�2(���Q���ַ�;����Յ<��+3���Y��mm���~�+�J̱8X���US�K��NeڪSv�r㝗u[��-��9������?l7>lA4֗��ʐ]������z��g+�%'M0Qcq�
L��U�lɃ�~�*g��Zfb�*�s�8����&��aj���[�#"&U��WDr=�p���LN�x�jB>����v��%��b±��R�	�Q��RK�}���������(KL�X�	b�o����f(����I�Z�3K�6PL�08ޚq�վ2L�"\����6S��0�M�ǳ;� I,lu}�8��<���#n�p��������1WL�/B5>_f�%�U˃�z��,ǟ�*�i 2��4��[��GޓC$_0�&���+���s�i q�
��C���,��mHJl��g/�X�P��|�瀊��s�4l�����X_���e\��*L"K��7�X|�M;�"�;tn1�E{�e��$�$����(F�Ŝ?{JŢ:��Pf����ѹ}U/Z���,dD)�Oʏ��%{G!_a�a�t\�j�:�uvR�Չ�Aۖ��8���$T���hr�����?��Kn��ZZײ�c�ǧP�][��X��i4,A�z�i�J�v�p��������SeD��vBc:3�����{i%  �&ڗI^H.l�x��<�XL>;�}>/O\�>��s��҉��Ko
�$����9_��?�� d��£M���6��4y�p�0���zl��c(��,�,����0�$�]s�I���	��,l+�Bt,w���5."Q���jg�� ��3�3s|�O'��;�E'��-H(A2�0��D��(2���G)urG�I�.�j\QN����������:��o���B�@G�=�Q�H��������#s�QR_L�N��3[͠�Ҿ�����(w�Hd$+9^��w��
��ܙu2.Pku��K1_���«�]!0b�ط-��lMZ%�Dn�q0Wk���Mˏ'��y�iOFz;�N�J���ۥ8�h���J1N�p�}M������{��A$H=��G��)*��d�U�m��]g�KY��ϩ�QF8y�昱=Ob!��n�M%1�n;� �כ���ʐԒ����;�W�Ro��ՙ"�a��+h^FY��:�D\�'XD�����F�L����%m�L�3�mb����,�����}��=��$��ܺ"���������l������ �鬸�!��������F�!�ׯy�mZ
���v���m���1c.���U]�.1fVM|'��mHٿ��½wM�������KꚶC�N]W�t���I�Dg騎|���j4����a�������������sJ��}��*���.��#���qi A��u��_�!�H0xar[񧼑e�����k�����'%�m~f2:C�Fp��T�zUd�"oB�^C�eU𫡓��q��/�;�۰窱wMO݁�P4�N��+��m�d���|E���q�Q}@��`7#��%���^�tΉP����.���:���M�A�}&���t�m���߾���I!��s	C�W�«�~�|:��Rxz;�<��\�h�=|R�SucIi��bjN�oum���H���`ҧ��I�y�ĳ��^t�.��x�*$<��|G(A���8c}A�h�΍��5H�k��sj�)US-���M���]w�xvC�d���30W`�-y����r�$�h ޼I��%�`��ΖHL��]\ Y_I����G<~{��jo9�ǹ?�_�.��	R9�%kP){���=ݨBAG泈�FZ^�ի�Q�61��*�}�#7'=M������w�*�C���	TQ|G7�f/ӝ.�T*�xp�˺cPh�b;���m�x�a�oL�sM�`�0��Oުga�`�&3'9���$�9��O'�Q�e)p�))��O�ɅH�5�
�<�B��	荦�iǞ����\�ќ���^��Z�Yb��J5�
�ʳ��K�h�٠Q��lU!��snD��H��T&�%�.r�,k��Y_]�.�˧g�K��H��ekM���)F��*s����*���o�EIy٭���-;1�:��߸�e���n�V%�Y�]/��l><���B8��>���[3�����wn),���v�vg�U�:}�~�\@���p6�x�C�Fy���1&�{εKٌ-��R/_(q������˜�p/��o�2k\г(����K��Pg��_>N0��=(W*��%9YFr{�|�8�JP
DL�Xqr#N,�O�h�Pa�`��e��0�B5���2�4��vͬL�>�t[�O	+�u�"5�L�ܚ�э�l� 2���F�aS���,�[� �~-,_����05�~qؖu���U�g�R�o`�$�2!qJOA���n�u���Ӷ�%rX�MU����;���z͒��!
�l�=����L��)W�U2��Bӷ(U(��X�[�t�����$-���� ��R������!vU�mX�ؖ�"kX:��E����~�qפ=n���ρ�q�O+�x�gs�w�4e�דTx�+� Bk���Oяn�K��A�=N��ؔ���r�>�-t�_�@��l�2+"�,H�(��)����I���"p��,~He}�z����Mx_��vy��g��K�\l�̥.ļ*!��~������ �/��R�&l�B�X�amf#	{�=�F�~��(T*�:g}8	[=�Ά�)T��N,Q�������)U��z��E�zc	�O�90����񼌄�m�ܞ�Ja�5��g���_��[��J��~�F�!$|�� d�b��S=΢�~��uP��g�zn+O}�G�k��f����a�.�P�Bm��G�m�qV��n�&��|�ԙAh�M�.s6}[n߀�O༟X�P�����NEA?�a�8�ȧQ�Z<,��G�
��"�U�����9����b��S�y��2v~ ��u�P��#Y��I4�f�lV�A��$o�8�Y�`O���h��h�9ߣ����3Z��m��b����k��a@g�\�<���7�ȚZ�0��#�5ML�l�7H�Hr'�3�h�ݣ38�6�|����q��u��m2=ޠEk��h𵊨º�8e��L`��1X�>�R�B�h�j���d'?PVK�g����|;��U��Va١�̰�#�]�y�b��,d��� ���~�x��2�{��k���:%�XnwT7�w�D������p�t�m�)
�X�
%	��]���ތ�3�Ldz��,�8uV�8p/JDͺs����RHÚ&[������z��{v�Z�̊�Nj���'�D�F=���w�չ��]��c�Gj�@�k��T2{��`��y:���f�.�$���T�ɞ�j>F.�_]�K���d�^du�s�� C0�i��@��)+�.E�C�y�^�x�("�S �p��X"FEd� ���	���¹�(�4�'C�� ���1X��(���Q'�����a��QL2:�����J}���@��Ǟ�S�;]�8tz:�;�,Q�2g㬂9-��� �K�y0����Ca,����i���uq�@��MXt�%��uss���<̊�����2��(#�!��U�}[~X�ߙ����U�?�SLϩh5؍��ſT���bl���X��dY��k�-�'[<Smx�a������@��`�X���p��Q��I��pQ��(؉��e�Ռ��E�|�{����4t�^��q�|������$�������ps��[�,Im�>�*�j����}S�̒s�A� �#�{u�	n!NO���Q��s/�N����|T�V_�	?��w��C����vq���"����7����ՠGa������	3�R����ot��O�;�UA�����>��Օ�m��u�`�᭖2��VV�T�d�ˍ�/�Wa t�S֚HQͺ��2��%,�Y��޹1-(L2-jO�k��� ���e|Z7p�l�%3u��L6��J��År��7@��r�TL�O��yDZO������ޣy�+�h2���oX�Z%I���#�H&��t����'��>TnP�E�"�.���u�҅����KR����?Ҟ�+�VL9U`Y���E?��Z�r�V:��/|O���X8@�� �O!�[B֗V�%JS����A�-��L��A~ɕ�v3 o2]��\8�Ch�#j��Y�:MC:�!�Km���Tl!Ã�_-�#�O��D�%�r�U�ZD�"X���zB�C3�������s���S_Ί�a�3�������a�R�X50�[�Q0��lh�lA�b�2d��ޞZWc��,	�K�Q��$g��Fȧ&�|A���3��p?�"��� t7\�8�ҲUY� �is�u��U�uhu��x����a���������߰Å+A=�\w��?=���}���T#���7<nN��R���d���x�Ľ�9EP���3�l���tbP���i�hoJv�V��Gkw�%��]^�d�t�чpk�����ݘ&���s��Z��ς����)�l81#Jw�s"~��d1�h�RM��=���O����D����"�"�>��Уun�윩���1����� �ղJ�Y`��Pj�]��`�t�IaI=�/�&��k���(&L2�/�f�J��C�;�����w��e���Nw.��z965�������H���R���l�~��� �U>��g�Q=ڋ�9����EJή�1~tֲO����73ʊ�J��1%�Oc��Ƿ���G���������1+�K����߁\4ڹ ��P��[��ή�F=��k�H1j��X��|9GQ*�o`k{��=׻�NenG=�>�Z��W�q�gM{cR�����<��!�U�(�`��ǉ4�c���%䓶���
?��6ȶ�s������bŚG�(������lox����a�11��-�]Idu#�k��~����Ct��O)�>�M�1��	��
�Mr���j��2�i�I_�$�",R���v�t������:�^(`+\��︠�V�d������-I���L������*i�ԬXdL�Wٵd�<*O�#0I]t����ҳ0�q�j���'�Z�/m������x�lhvK��I䮐ל��|r�z���.TޙQ.[�/���"��p�A�S�f���5�La,"���SL}n9}��o�j0�o5EɌ`b�����p����;�Ѫvh������H��	0J��f5�.��Q(y}�>q�J�zy�����6���jC����彞J�X�XG��M�(���O_ ��:���x�T/"���ȖB�(r��o�֤M7�:�6T�H�Sܚ,���,#�:g��:�n�r��1�|M�SR�A�(U���Ϣ �2���9�J��w;H��~���Ԙ��ۥ&w��i� ���nYS�k8#�K~M�-�+pL����t���Ӱ�N]u�g��_n����֒�*�f%b�?oY�ܩ�A�>n�k��Mc"��A�h� P�e{��3�&j��v43��c)ȫĵ=��Kjf��������]juRI����R�9�/֢q��5��2�%�� �H�A/�b
A���!�o�(�'�h5Y%$�|D�Q�D:<Y��A�bZ8���9�1��6�Ub�x���
y�5!� &�Z�
Y8��d)�)�j܀���,|�2ϖ�@���=���Z}/r����Q��\�+=ND�O:]Ё`�u�.ԭ���ͩ�<��Rk�I���̹�My�J� �hU��Cj(P�Ij]J�Y���D��N~7���a-��.�e����'��v�@Y��us"$QX�l-���)5T��Ȟ���H1:�b���f���zج�"�D�].������~V�s�E�2G��",0=f�3�ΌA��*��$�7
�* ���w�?�Ñ[���R�PӬ�=���.��G	DH�N;:Xg�g��D5\��Q��f��ħؚr�t0KҊ��C�,֥Q",
Ne��b^�+PnOoI �������X�����R
����O�-�8>Q,���r�5�=��/��:'Ⱥ������dt�=�+��IZ䅵�7�q��^��>Y"ȟ�5	w�!Ru)��@��h�R�cV�J��	jzP�,��}�0VrAޱ����¢�����@Nf���>2i�� x2��>����8�f�8.���jd��g�`u�
�)n�|��(
ƫ�	�O���(�&��]��2vv��\S�H������5���H׊��7݃���݀D�4k-ձ��l�%�т݉5�P��4�o�xv�e&0%�rjQQ-'�QI��o���5cx�����s߻���1$��戔7��=T~��V�� ?8��i'�����8&����$/n#i��g�7n%���;J���_�m*\�c_<,��X�%�T�1?��M��:����p���L�7����[�� �)����Qq����"�ɸ�J���hH���9�P@<&�D�[��"�.9�4y�̉�7���	I���"���OV�Q�[�}��1d��r5�Q��m���os%�)N{�7{^�vv�u.��`LS ��k���VmR:��׎���:�!YBuU}��g. R��j �v_�-��'�	b��!vV�t�gW�Yq}�$u�8t6F�C���7��z9S](�m����f/7/��-c�ɼ�ڜ�L\�c�t2���f ����LS��LV�,��B��3��[�����]2��P�i��-mK}F����d#}�
��w��rL$(h��o��h�a��8�������+�(��=����s�~�|?�s��^uk��A���	ؾ=�J��9t.|��`�%���+ ��ߗ���E�^��������S��X�����p���?��Z�ӰĆ��y�2<)Cb�;e�1�k7�-���mx���p*l���H�r��<A`
�39X��[�pp�1�����F�G8��ei�IK�%.,Ӌ2)�`�7�9�#��l2@umqy	ן|�OuA�/��9�d�+�A��@C�4o0����Gw��ь\HI'���"���q]�r���o_��6��9VƱQX����[���J'��d�t���V�υ����mA���.����ʗ���^KTGv���[��+�	�ZП�X.�6a��Y�ͩ����,|�"��yK4����9��z��矆�e��;�� Y�D�G���S	`��R�q���Ǧ-���g�Q�]�J����J�B�ڪ�Ο1{dP�5�B�` 0���JT������:�������R�@��gY�H��2g8ZҚ��ǡ��dk��E?V�zX��������8®�e*�pa8�zE}Rs��1��Lғt�(^�p��x�wܱ�Ɲ�>��hY�P[��`q5�z��D �A�Ӑ��nA��;L�hc)�"�ҡ�`g�V~��o;6?[� �-��uNP��cOB/�6x+�H	p�R�r�����p��;Yg��oj)�/3����^���h��V����s���ʥŰ�x���m�@�qBܗ۳��֕\{��:!��j���<�O=��+̘�&�m�/���o_w=Qk��Ze���}�A��,�Ik�5Ȕ�Ԉ�C��_@E]��w�ZCyz]=��L<*?�6��2�<Ճ���"5�D����
UYs����a?E�Cl�I�@'Rm|��,15~�zF\pV�)����ηz�[�ۭa�k��e 
&azb�g�`\�JK���X7OV��_�{����<|���\]�u�c���|q�P2���V�kZ*V
Q���HE��%
1S��u�ӈJ7�\�N����8f d�;�MK��Ʈ�u��Z���@<��Y<���3z�.�Hǵ���$Y\6G���	`�ɍz|�as�wr�����;�	"U�'6�sʅ�NGO��5;o�V
�\�'�.C��ZT����~�-@��EP9���t�"�԰X�yK[��/�W8�R}���pBy��%��i%!�D^g��ݲ���߆V���1W��GTLd5���`�g�������h=��!3������0���Ұ�Y���1����C�Ԕ�Nq�����T�.r�Es~�LMT&��j�^��n��<�i3��!Gq"�^�@����S��`"�q�/'g-H֐��.��=)�%�7x�M�(	�X��#b��N��;ec- �#�ƁN3HcIc:5�Լ�T-$C��(�܋ɢ	�ԅ<��`}I��1����)C�pb�TKh[��O"�0,������9�{L�c��><�Z����\���=WbD��J)دԁ���0���5�� ~`��Iu�����#�UR�M�G�U����U�E���D���XdvE,+��z,�݁�����@��#��{��1�;V��e�P�@��g�T�"�U#]�ux�2�˟ݖ���|��'���"��IY�"��٪B�7/ M��t2��V|��-	'�vN�9��}���@���Ȕ:σuh/�|���w���)�~�`D����Y�:N=�)@��@됌�c{�D��GAB߳��ݲi�⚆2�ӭ���U�4���u�r����޻}�g<�\��[��{.W뜌v�]D�-*��l�L�*i>���F.����:6e׻�R�}l
3!d3JaF$_�Or���诏d�`��&{��:����&���g�֌�?^��]�0�if"k��($@��'�k�_��{ 6��a�~����.C/�ly�L�|����gKU��q�hSR�!�m����_��>=��#RR�7�5����t� �����Qs�L�D�ph�+=����ɯ�jC'c<�;ο��jnC|�q���.�_�m�L#cA�Vp�\�B�#�<��Z�`�^ԣ��3L٫��^D+-WUa�{����vd~a_ �z_��j�(Pr�H����ua�V%�_��0p^�e�!]R�<� �h72ޤa^�;�Z�5���2�Gxa��,�{���_�%��
��ʞ�^b��]J���B,�����O��l7��U��S��s�(�)����Y�:��5pS>b��|}��M�Z2�z�Z9M.���}n��k9h�S.�M���HW�q�[����=�}M
D�*]��tE�M>Ǫ�Jr5@�ʖNFJ��T�.�4�� ��x�xz��۸�|L��%O$��=��tZ���/���XP�&cu�l�qЉ��z����Љg_�^�Z|Կ)s�V�pR�Ǩ̻��ͷav�=����ֶk�;�?ܖ
l�=�)D�
8��Lؚ���9�.��Ըt��+��ЅS*��Ft���I�T_H묚ˀ����#������;�y�����Qg�4��sE�Fb9x�9�o��Ƅ�Y\�Z:I<Pg��n���Q���Rqͻ
	�|楄N(C*�0�c������1Ǎ��[}{�*��s�W�}ZWOȉ�W.���D����/ L}S]q]x/�D��{�9��=��V3�'.kO����W��1��)w�_8�yK��j�Ô�݃r�[�ێ]�QZ�"�
4��p��;c��TNXYq��2�=^�ZБ �S-a|�ֹ	�4r�lM�umi=ʏfi�t�_��p��><gB2 �4X�b<��"�m��-c_�â��y`�~�;�}z��Z�'`B٣`��Acs��zF|�N�O���X�?ϗ�b��P���<���DQ�?�f������`�?�ϒ�����qp�ɿ�NJ����y���纔9u	��g6W]�S�9ƞ�`����񟦏�
/��rxk�6��D۪�C�:��o����X4��=<��~5X�1UJH�s�p���?���`?��+G��Q��*�7���X���Ê֨���������F�r��ƇH!Lv�%=n�i�M�r��d�"���N8`t���`Os�9b�=1Z�ج˸��
�a���U��%�Ɠ�rC�I������l���oȫ9l���c�8����N���ђ�{V�cj��E�_��^��翘m���6&�qt����k)�qX����P�����S�W,Z�gKR�oFp���R���	�>��}�&��A��R�ޝ-�Ie@�O�`M�s����\����E1���a�l������~�Ŷ�����E�򬮒S����!:�	���xj��ւ�Iט���0fm?N�Ӫ.Ǵ��ɦ/Msh�|{x
�u�$����!�0|���<;�䠘1���=`q��P8�W6���p�tE��w��g�F�"s<�I�}�ci������ ���?�sP,��|)��Y��M4�Sae�u�h �e������F�~��X|ΖUQ.�W�����ej���O��:5ؒ�C^��bo�B��
��Sb;[�������K���g�@�Ðe��G�ڀt@^�J�f��[$��]���y+�`��Bº�:�QE��B�˚e9|�3QL����+�«�BUZ�9�vL��@�`y�w�F����CO��wx��p����0JP����U��BDVo��]r��
`~��2?���D������*�� �ߜ��3[��Qd՞�,�h,C\Z|�T��7w"��������}.��)��V�1q9֠Hu�#A'��#\F�tZ���b�/Ag�j� nW�0�ZF-��S��I^L���u�E��,2)r�B�^�f����X�c�g��JA=�������E��d�g��׋�!���,h���;�|��_-�r^H��SS�x��v�{̤�=�c����ǽAj�#��Ӥя���c�N8����Ƕ�Lg�~��<���`5�n|H��	�<��D�W�{�vK���R҄A��Y��-���a؆t��L3�+�V�gq��i�Z�u9�$���d2�(��|\㿑ݛ�Aq&��0PF�>.�e�e��b�-�=S��?*B$x�,�]x��p߯������'j��-
�7���)���?��WZ�p`���u���j�N��E�~>��ц����9'�ݝ��٦j"�8��9�Ѭ����[d��=rk�*'�*����4FL������TL�=���56q�>fl�7������g�ȳ�^w.~��=�*�S'�3O;��~�kZ������%�+�o��?m�!m�T4Dö��M�O2��8� �4��a�~�ZDk5�⋜�`3@ND3!N��9�ru�Źr+�D5=��٠��[����ڴ���Z7[�x�\u��\ظ�X�[��+���D��?��3��j}P&l�T��
=e�*�@��Q�&�ҋ�K�f�2��5ߒ�!^C��Wj3�m��tE%3�+v��)����C`�JI�
����B��/��r��n�����XF�|T����.k^(����F�p�Q��RJ���U#b��m��f
o�'|J���e�|�°ٞ������[���K{��H�d���=D���g5_9y�Zh��^���K_!�-.?-+��C3:q�?��\���� �*j?+�/���Kr��:����I�N���֮������T�Tɨ���Yk�B{�1HA�|�Y�����:!�����[��&Qw
�vR�ԥS�P�:ƒ+uk�hm�z��%������:q�`Dj�<��G's�W���DG�x�� ��i �o<�{.��7��[iMM�Y�	.�5�`��3��cA����r�^z���Xg؏q�G���cEe��n�kd F��FA��R.�if�r���z��s��������=�w����Q��.���<;Q���3f�>��RQ�b�'\F�4l����j6�~�HSgx�l[9:`H#�]5�W�+��^q�6Q|�ۄ���_�}N��%�Ǎ ��S^5
��}�w�����)ƕF3rm�]�)6]*��M�ܲ'�3�E�Z��r�!h�Z����+�_`��%a9��w'����E��a6�A<xL,��km�NG^��u�5����׸��ӂ��bP��91����s%Y���b&M�f$8���L������齎���:?����J^��~��y������]٥2� ��Us	�q���W�a��L�۫ p���m~��;�]�HcUz.Bs.���L��#�o 'b��N�&n�ϼ�^q�Y�dc�����ӀJ�W-_b���B&���YF#@aR�P3(
��4�r��C����?�7m�~��ǲ#�����h��M�t��C2m����%�,��9h=	���fu���l���@��<?��C�3|�`����i�OfY*� ��e|%�YƳLmIbmm���C��bvב���k��`E��<?�E� 9X���RJ!(��~���3s�*<:��ւ6b�V[Q��,4o�P�Y���N/�I�����1�\��c]���j�A�A8*z��^#f޽nJ0,[/9ٮ��UK8��-;���J��{I�ϋ�=9Iǆ5��3�`'`��6F���C\�kWqɹ� �?XCk����0��(���HW�.���Q�w�n�9�=�*�ن`>?V�:��~v�@���i�C�;��x%���Nx\�G��Xz�S������ݍ��K��6��ڐ����cAc5��r�O3]on���b!Έs}����S�k�9q����*���,�2��Y�`V�����n�FWR�3W�}c�Pe�DK05Q}�){&_�uH	� ��c�����b�>d&��7i��ާ+�(԰��{�U2�Dqt��&ލ�+MI9;�/F�3�Z(0��SZ=���d�m��+T&/�/[N�nE�xP��!�w��H�i
��˱���q�a0X>����v�"�4������J̧�!�7N�Xʅ��и�e�����աSU���R������
A�h{����D"�*�3�5�N���X�K�ݥa*b��ݱ�9��~�T~H%+:����KD	�!
�ޚd���p�����$扳�̽��̙y.�� 6h���d�ل����SZټ���Ŗ�$G4�ns�(�~<�������>E�f͡����R3���d%�������HR�K]��N΍��"�e����W)�7>�\q��U)�%�W�O@�/l��U�.T>��f(˸��;��~�CU�-�k\b\r�L�U
�/@?1P�jN��G����.��X��O�<�K2`%uc�|����(���/�����s�Z��m�Jℯ���]LP�S�p����3��J�-�rD.�����1cwCW���T����g2�G`	���Eb��y'dd��s�@���(�cnN4�7+@�xg��%�7h��jK�M-Z�*v'�����t��чHl�rњP�ybu�kz���=���k�Զ�ǟ=Ni�s���C���ޫɗL1����k ���5��x��n�|�+�r�[N������l�n�s����D5��(Ye=-L+�1�{���G�tm&lY̑/e��]I)
y!6`yc!X���:���,�x�H�-^����rl�����G�T�{�*]��O(������?No��{�;o��J	��t;�B�O�])�G�Ԍ�	Ё
THq�j���xP��Kd.}����Gd��G��. ����joBo
�_W�������~ƍ����KT�4�����2��r�R�F�;�M�	O������O���B��-�H���tQϬ�Jz�p�m�a:f�Y��?�x���LU:mX�,9T���֌�G2v�^2��4�A%��mO_�k�=-�>w;����9�vP>� �Ծ`'.� ��lܜrpAV��G��� ��3��BOUƪ��#-�pH>��Lӹ� ��wZ��,Ŭ�X�qr�٥�EY�!�����i(�z0w:�s��y�6����?���JO���L�W}�$whU�/s�Q�L���r� ���uu!S+��*��f��{����0P���-��ed�G��3�m�=gM_,�!���q�I�G�ݯAy�ݎ%0�x���2�9¸硑T�TSdV.�U*8N��++�?������Ƈ^����>�ZK*V(�[3G�ʉ�(��(T�.{9s�58��m:�zhR�2�K���x��[d��,YƷ�՝ �)����p�R�P]�S���B��c���O1���䖦q�#J�����Ti�3�?�Ӏ	�*�Z��&db�Å?�>��Q��ᡋ��mI������\�G �aW9�1�T���S�!,!��غ�fp���.�"&G�b�"L��ݯuڡG�bI9�G\bl�J��X�K�B�N��9����b��S�/
y�3�^���!���)�/�jx����r��U�4��� �q�^����S�ЩAۦEף��Ѳߗ%;�f�Q���`���)NX0�l1�[�D]N��w7`L��y��'��M�i;�b����FW���(�Hف�J4h�9�I*i0��>�����ټDvPW�6�>�����H�cOӸ�SK�Q�6X���RG9�����^��[�-�lF��tF���aE����`�=�sQ��[�5e�]�P"i���	�L۝rN��7�O�	E׹��mT�c�E�~�j#o����Mp+�R�d��F���.��R��7'g)?��^�u���K�Q�/�"^^�O�)@�u��5��v�>%�^��b(�М謳���o�ݔ�s��.�D�qV���G+on;l��Դ�aR47�2�>��P(�S;"�ڄ��@����)\4A�0���i-<.ܶ��/0�ݷ�a/�궕��ߛ,bg� �����5�)Aߒi��Y{rܪ��XF�}��O��J ���l� Y/�;���}�ۡ�J�{���%����v�qY͘Ϡ����z䩺�wpK��ˠj�Ç��*9�L���Ϸe�/�h[c1�5E�Eƌ��Бz>"�|�i̡s+���m�� �61h����s��M0K������������VAPrq�o�$3��	Ց� FE���N�^,��1�����/Ǳ~�˕W�s��D{�j��ӝ4LO��j-�r嵊m���fS1%�(M������ɣ�̔6>�]�b���b�d�/��aQ�����u��g5q��u{��B�N]h�2J�� �����#� �J�%���~A�]���5wX����^��\�Eq�ʊ���N�����;�+�(���Z��g%ʺ<>2�!�lh:�&ˇ=��\����Vx�jj��s�������l1�?�Eހf�D��� �����00���@�6ُ�\}.ewUao��(L�}Lb�^N)�3͕�N9�@s�*:B����M�A�Vd�RA��uˀN��0n3XY�}a̹��N���SÀ��~�ְ�(����-�w�<l� YΟ�0�]/"
J��qE8֋d�K��y{�w��1A�M��^nh�>n8fB�>nL��{�k�D.�`E�oVO?�֒}����䴛�lP�Y�݈q�������<�s1��is`��'�q/!3aSő`��ʣ>��q	��B�o��2�?k{z�7E�L!�k�j�	��<�0���og!���������M����w���G�����M;�0B���hAyF���>M��n�Zu7W&N|K!�;:w��x�j 8X"�����S�^�$�����m�0?I�B��h)"��m7���`�uAM�s�s���@=ŢMCF�����κ�L��Y����������kU�H��5
��g���D0��#�%W�J�!�|�4cP�E^�
<"���:��M�p��#6������&.���\p5Z�S�^G�l��K���s�Ŕ�����%�z6ue��[{Ѣ
��J��)�PJ�G�Ժ��S(���p�h���� �0���{��T�t�h�f뜶m�Ǝb���!����M��<A����Q��j��g<`oo���`?1���1�q���l�p�䏻L�8�k��f�BH��\��ڪ��\�$9b6�Qeog�nm����0𧼌��� �1Rc���e�����<d
:�{��:��B���f�*�w�L�J?6�K���{�x}D��w��t��7�Y��^�/���z��$VcXY��o�+�X8�:?�����i�g)Y��Ñ�V8;�c��-��؜]���QQtߊ�j,���D��a~b59���L����CgI�B$0(!�Z<�k�;�)�RRE��(��}���pRP��b�^����e����	)�QaVvgX]fRM��u�+���T3H|ѕԄ���O�����`�}<b6:4�6���"�5z���S����/��IJ2ZY���
��(&Y�#�﨟G��í�Ǻy�O�`)�HP��7�)��Q�H��a{�g3f�� ӈ7�k�Tq�Dٌ*�>GZ �.>��Q�(�xU������$Q�8����fh�z�ă~�ͽ�G �B����Ιa���<��&��J��]e����M�avӛQ^�� �Dp	�ݴ��\�ѣg�rm��Й	���P@�^i
r_ϒJ���b�$Kj��j*�楸���W\�:М	4�����B��b��g:ꚝ#G���l$˕�����6���<j�>����:���(I��Z5�T7uuJ�7嘽�V�K�QP��r�X��1M�M�����\{�cWp��a@W�"�"��)�Ǘ�-_rB}��8eM�I���y1��k�>iy�E��t���H�b�닋��q��RhF�l���0IB+�M�ح�'���e��#��=C}g���'���ب�#��s{�& �L?I\���q`�p�v6��7�#�hܮ$ ;��21����B��6����ֳk����)򋄻+iw]}��V���$Z@$��i�F2�;Z�����g���~t��uHq<��y6�]��:Sv��v�S�0�N����2w�^,�<���/ȼ�"�ir��u!A��Dv�����l�ƙ��I_�\���V�A�����/�${>:&9�sϲԭ:Os�O�ji�6މ6��ßcJ�dBOEa��x3�R,�	Lj%aK����-��|o�
vi��k����G�������|Z���dX�K���ڢO�!Ad���A`}��"9\S}�]Lڌ�=��t�
�"f@��N/�I�r�`7�5���B$��\p�F����6$��2_�.í1QRk�n�9�P�����-r�n�xi�G�=12Li�.��*��_����JM<����� �&G!�oU�N��RsN� ���3�����W�m#
���]Y ��O�ɴ2�?�R]�!m�.�0狊����&TT��T��7����y�c�(��3%JD;�s��~�pVm:kY�чs�ib�?�P�a�d�I�6%���c�S6�~+�5R!m�����e$�	�m��� n�z�~���n�s/�}S���,q}�^�=��/m�g���T� �����<�ЯDL���^6[H���ʦ���x�N����9���m}��	�����s>��G�.���E�#]�_E(��p�H�^��'����F��~(̶D@�7uv${���8y/�о��Y��R]k6�J��[����ϳ�Vʒ�6V�4�8�(����XE���f0�?B�,U�P&9����g~D�K���d��}^7�z[�O��ma���AHc�!��c,g�B�?>J�����(�̥�/�Q�����<���=�c`�D������_���>�qvB���WwmAԹ5�;Q�IS H�C^���S��Ȼ7oI�3�w�0�2��^^�<��;�nMϊ�?����y/��V:�ܓQ/��ud�b|�����l���w#�ʑ��es����+���wĔ�V-����5��2r��&�8湁"��̮�p����X糚1�}y~������T���&�E� ��LU�!����!�mc��v!H Q�/�P��F8��ڋLs���aY��\P��:f0х�r��E	y�r���l��z�@hXb�� �	Rq�񬸙AΈb��?��	ӛ����0}돪���~#���b���=������ݑ5n�fͱM<{Z���|U�zǓ��4Q��'w>6E�RC��M�#�^���M�ͅ��o>*6�{�h#�\%���L�g6�6OY�?�z,y�A1���g���%�o�>;e����tiD�v��i����K��ƴr�Ũ¼kG5�h,��K�~�l���ׅ�D���]�T�.Z��wח�C��T��� ��H
������F ��6N$���'�c�a!Vak!{e�Q�����]Aa���9P"X�k�~d)��<�)�P�ׄ�����n�F��=�8�".0�L��B��b%6����:m3T��Gt�����o�5��A��eG�wo����eQa�R8���Y2P��3d�q|�j�$�*��tz{�"��0�x1�f<�I��#
Kء��&`O���n3��M��E�4E7�'�?���gFS��Ș�Ir��ʀ��yfr��D�0 ��nE�JTȊW�o�+��#��G���*�xq����&�A\����I�7��	y��� X��/��c��r$�)�{-ԱjÐ#c�1p�Cj��5�Ubv�H�q(�{(t1E
�@Ŭ����$�ο.�a��mb�R��f1� ���>A5o�)\/���F�1[� qI˘,p#i�>����$�wJ�_�ڽ�s�_V�ϳ����EyX�4�|�r�Z�c#p��Lp���S��q�Ԅ_6/ V��i�)6�q�Ꞓ?���%�I�]?�ho���l'�f3�-Vz|�����������g;� �R&K�U���L�1T�UH��Q����t������צɳM.�;$�i����`?�:�ǲpcĆl���)�f���ȭ�}�e�v�E)�$"߸�sb�����p�^x��*�b�oi�_,�o7�&��U4<�/P+�P�x�o�LP1�e�;l��A�gٗ:���ǩH_;���V�L��_zh���!��%mZ,>�wL2�чV)���;n˩�S�
k�&A؉�?}��'�o%~U�<�,��b���وU8��`�^o	�d-%����C����f���FY�L�;]�t*�X�o-�_��w����6 �����ފ�>N�_��c����f���RAe1Ѕ�7���1��Q�(���D����(i{� (���p�d� �Q��0��q^"=�4GZm##�3�	4k�eNN1���Dʆ�iqd��nNѐ��T�(��`Qs�w�s�r��EC��=�ݻU��*!�m��=SI��������.Nq.�Q�A�	b��@a��>Ѫ3l���z��?��CD������̗�I-.;垍�	���7�{��U�p��ٔ�]��K�,A�Z?T�����-zg���:��&lB��4��T�<���2[�QX�6T�8=�<pb���3��O
Q�A�3��FϾ� / ������ӄ_�(q2�56�X��i�Ĳ��[�3���N5rq�l暃6�r�hQ�>���v�o�;���������4���<��G�0PV�#�·P�I�61:goC�q��.K�yY�+k��7=�`j��#?�Ж[���Q��\ϴ���SV������Ľ��Q@m��8�q$��o�d�~�ރ�R�-�LeZ5/S���,���k:�H�}��������8?��K�����H��tN��DY�V��	Q�1����P6Ys��p�E�U�|�չ����</�PK�j�����W$0��nM����f��w!GB���=Y"A��۹ �t����U%[��-fo����o�=���B[S�.�utE�Z�W[�$q�5`y�L�d�=X�Q�v����X���b�8�^����\���%�9��͙����؎Py�D��Z~w�9
�gA]ϬHP��h�_h�o��b��i{D_� #@.���	�3�Xr`� _&�S��NS�er'�:s���[��(�� gF��e|��s^���"���A��+>�,z_��1*����&X7��0�
�ٓ
#���@�b��
�n��@���(�HR��~�g�y@]8�K��a#ڮt{.L^A��H�K�S��}�-�#�!i�\񯳯WZ*�1��]�&��J�ђ&���֝Y�hm}�h)��S�
�U���9d���1-AEB)f`u�6�4�기��h"�t�5"�X��'h�>Ig�G�k+�G�K����󆤰�T�N��&@ ���=��i-�W�� }u]Ю�'j1�p����i8D�\��g�V�����Ev���@3�'~��|���b����-\�ofS1=N&["M�z �6��Ƈ�4��wT'D ���=�B���c������Lq`�b��{������ О.�j��K�Xo��&�K�پBж`�g{���B�&��>9�{±=RO[�@�P��y"��},���?���;/�$9� h��sѠ�m��L� �J3�42�/�t�1y��� �d^����G����nu^h����U�JX�t��;���Qp%�m��Z:i��-'��j/&�f��!��`������5ê��E�9qޏ��f}�����(E'���� ���řHM�J˿��~W.����i�+��r?�����gCj��oXa�#��/k����4��Y*���Hg6�Z����s�$�����d�x�kj� �z ��^@┆�3)���4}���'����I���-�ԫ��ً,�p���~M*�VNtV��I����t���p&shPW.��%�WGHt�y�����l�p5�0y^�Xv�N��s�����^�����}�����/%����L ~ ��9��	w���< j ~M/fE�,�Dg�韪�����좖�
~�d!X%�1��n��P"5��.*ޑ}�soK4?�t���U3 ʰo�p0�Z��<��"f�V���R������n��@d���ջ3���*�k�n�wJ�e0k�{l10D��'�&��`�z�~��S��0����i4^L(Q�>��~�H�W��UD;�HT�W�#���40b�7�&�JG�s�H�����x1B�r��~]�TN�����?�j�j!���snMd\@d��k�zR���W�.~��3�~���f	x�2D�+��}'Sv�S��ˉ���n�dsjM�܆e���m�EC5�=�S�~]�n��Jn5�:w1D �ן�i��`��`Y�`����*�/�:JxI'���N�LH�ϯ�����l!ä���W���?(��h���m��|��/}��5
�[jrӹ�t��ȣ,L{��B�� �妅�������h�@KF�Z�/144c�y�r����m!���`lG�b@|��[�4�ݰ1^�ɫ���X�f'`Auo{�UC­fj�[ʡ����zEMg�1]��.D��q��%��9��?s��˵�'1]���v�r��(������H�1G�>�?K-L�:�@�EI�نe����OF7mV5}�C���� ���m�#��F޲���J���������x�_#�2����4ݺ
��6���OܵP���Z�D��o��&gϣufg����� uEKfg��a��|��F�龝o��r�Ѽ@�j���X+���eA�w�}���@A�������Y)�h)$F�Ҽ�9�V3�gf_ώݻ,9ql�v��y���Vq�6���v�����
>���m^e����
Wpc�ʶ��\��	�t��t�QE&-	H8��K��kj�A�A�6�
:�i�~ ��d�P�~��c)XK��,�r��C�놶����$"�W����%�\ׁ|�"Ɋn�hgp�a��|��,�MM[6B��	�Z��Vyn]�]�^���"�@�0��~�
1g?~\=�`$<�P��P�%�@����f}Н|���7WU�д����K�\�����z1h���lvͺ|nY����U��q���]��8'g_����]Ŏ2�h�O�v`�>p�f�F�S=�M��	�OҦ9���lBn�JӁ+:� �Z��~�H�kRH�o�S�?C�P�`����A�J{�d�޿t�\U�?�}����ٮqܽ]�Ef�2
���@Jʸy~Ѳ�!� ����"���o������*��s-�7O��t��W��Og����]^�n�J�Ȥ.����S^k�O��+ɀ�Ԉj<�>�MB�t��㋬�e[��k���p��e^����I��J^S},��3�Dl�>[�u��W�D��Oo���8��/�^J�{�"�ᜨ��-!ww����R�ˈ]Ƒf&/߿1�&<����\:�d�TД���!��⨮A�Uw5�D�L�bh��IPg��b+��K#��E�%�s����Ft�~`�(���>��E��ڸ[�N��(���3�����Z�h��?����	p�}ו�u:j<|�2�ӥ��Jyx��LT�72mZJ�%sR:H��<�n݈Ý�ʴ�%��D5�je��p��aZ���<R���fC.
�ʙ =p�2VC�R�A���d�C�R�N_l�ۈ>�xA�R����\�
�� ���&U�WND��yv��:�Wm��ZS؂��rz�̬���-���'����ܥyʘz�ёX�!5䟂9����S+���@l��~_B��{R^������}"�fk� y��Ds��!n5�I(���$V:�]؇X��fS�0�󕜚��c j۠>����<�9��:B-g��%6�Kє�ȰqyԽ����ֻ�5�ib|�|����v����
��mb�y�� i��Ț&~�cvmo$��q,I ;�o�,�7�Փ���f�����s�ryɇz��PM�E�7:pdc%9�"zY��A�'��3O/�`���A����@ј3����u]��E������-ݛ�c_���:q(*G��<��,bUݾ��-柇Gzpءe#�3.��:hF�� }�F.%��$��,b@�|���T?,AR���A����(��4��,�=��:��5�=��5�g�2CZ���#��R
�b�ѧQ�+�������v} yl��<?kBp�+E3��*�W8+D�����!��p?/����.���s�`VĲE����Z����t�3�}!yf���duc(��b���ytr�I�ɕ��9�*c��2�x��v�	ޖ7�=Od�_���#�U�>�R��##2圚/�+=��j?�s"��F���7�}��)�曲��_�!�s��сp��*T�?�j���TC�,�2�n[	��g�.���£X�̓�:%i�s��o�6��?O��Sg�zT��<��R��+%.K�;8g�l�"�_���G���3���b���8�a�X��xJo���p_���:T)7uʄ�Ό_Mdv�M[�N;��Xz��f��I�����f}
Л�KLV�o��ߊB�#̲-��:�ʆ|HIe��쳄�h�Z�&���';9���9G�D2[�nۄ;����=R��#d���źt����`"2*�V�䝉�/�,`����x���1����o���gM�ޡ؇��5�2r�zר�1ٻ�n� �K�&p�beڱ���^�_e5�q�H��ւV�ۿO#Ιg]j��'.�G�H�])��SdE�Z��`�����j9�}���[����v)d�&�N1� ���.�t�'���j9���P�K�ph�tNj�����U�PBu�ԃ�P�2f��<j��{+d���#1 �e��,�
EV�����U�b�nT=�}�p����#�̛��khT�7�;V��XyJ=�Z��9`d��F|�@]: Φ �(�-}2L�L�=�2*_B5>.�)y�1e��<�4g}�I���fP ����^Ƀ@+�\fq�{9z����A�J-�����L�0�m��~�j��jt�
���� �!�C�K��nX��JXeo��?����?^�%�~G)�)���X�
;�X<8��2(Tk�q�Un%D4r-�s��<�I��9��u�-,�V�- �ӄW�o���1�d���r����E�#���~�����i�~�$M�S�W����T�y[.�����!>\t��$�H�H��+�o�AlKi���	�B\�b׀��g�c6#�'��j�J�u���Z�S��p�|�{�>�0���(��?��A)ޑݥR\5z�;7��f8�?�f�v��I2�]�%?�8�E���l�܀���7��z�Y�\ŵ�y���>]��.K�7=�dǳ��ͥ�,�� �������d[i|��%�y�dĬ\'z����j�Os�N��6�J����E���M�0R�v�� ��"hDE�x������9�>��N�Ђu ��f�6��AoL����e28�%a��7՜倡�ⳂWH�T'��BfM��4�d_T+�5��D�������dI�V�n�>W�����)�|�OBV���s��J�5���^�`;Ȅx� ���gN��%�C�E�95rWw����A{�BŤ3�"�EF�j#��4�("�����c�}S� P#oe�Oa7�{<j>Sf�u��)>��E��&ڃq�fƅ<��������j�E�S��2���~�P�f�(�I z�Qp�!u[P#O�ƙ���~\_,��HJ5�[�W�l2��*�/��FFx�1O؏\��a��M�|LN<��_�:���S��[E����qb#��q#�\�=�>M"j���3ؚz+AXx�7yea�� B��~�'���_������GI�j!�����a�L����r�>��t���E�jN|Q�#L���P��<���j�L�������� �*�T���B�S7�̻ �n�k"ǰt��:udP��`�������f�$Ĺ:�2sl���͚so�^Px�h�_�}3�#�ǫl.�++�`���2�&ۉ�a��
u
�Ns�y1�Q��q�HZo��O�2���K�bWQP�w�~�	t�(�EB@*7i1yE��-\$X�դ���@v��U�r�xgzW��u6�&_
�n{�W�#�����d`�/��-�p������F���M:�l��{Z�;�M�����J T��FE�L�+u���$�01�Dl&�hJ���ٻm'��
�ڔ<f��z$lm�%J^�
������#ZI�$渒���� ��M~v�GZ8�c��O��J��Nq��@@T���B���/���?.���]J�o!��b�ɣ:���qq�Lb���"N`�fKA�j��~�Q��c��\���T�RR�l�~+ֿ��5Ƙ
u��!�#��i��
���� ʏ1�qT51&X�y̌`��.���	q��v�i��g�/�@�|���U�"����C#�{�U�1�r7dW�M�+p�h��U�#e��S������e����Qq3����X��n+H�)��[x��V�%���������'�����p��P����'y�V��#�r�Q]����#>��hČ8z�g�n��=�wO�C�2�5
�d#;ǒnʻ9�h-���O�; =���V���Z��s�I��Y/��-)&�t]i�Xd}��H81㒪b�?�x`%c9�T����B����A�3%�2!���.+K��;4��������*�0����H�u]�8t9I�n>q�T�� �{(���:@hW��+��n��қ|-;��k!�{���]=�區+c�⢊���]W8"���_�B5�JY����������Ȑ�����F�_f}),�|�a����B�bS-щ6H4��D�QU�B��c#���z#�'��א��=��|h7�~Ö`��Qaj*!�l�{��:m�YH��wV��)�jYH����T�Ӝ�!*S��R�s!�L8��߂�ɾ���'褪ɒaUH�*Vk��M�qMpmպi�EN�W�e�`���kR��������|U��Ņ�K�d�X	�lB����6UR�>��ydk�I��FUS��檷a���=�)�K�Η���3��}9V�����/k��3(  
�D�������tQ���9z���#~��ب�^�����-I�e<&d�N�2��N���D�L>*Q��X`X퐥��?Z�|{�iT��n#k�v�� �}�v3�Z!���"r�ΉX�L���(9Qs-��<4���9{�y����p�*%$;&m�����IT���l�	�����´:s��Y-4���T�_G��gX ��x��L�(N�wߖ��N:u�9�}��&L��~��:��#I�UK3���8�z�gv�s��>�9_���O�/{�;�4�$����������^:*��{�vo�o���(m}Ӫo�{�/�\m��x�p��6��.,U|O{z�QVF� ��4y��Xj<�g�u��5]�D�&�>�\n�`��P��dR��54v��jL=�~*=��:H�	�J�R��Vn���� ��r#�.Ҽq'G�-LY�r �f�qD����^�U��&��T�{��`��Nil����WY�k����A�����/�p����
�ú��G7�սm�����b�̼����}�pݲ+�����Zͮ�O�6�#g��<�6�:s����D���D8IV	�j6țR1���yp]&�6��-��"I'���"��b�H�$�>���S�ڹ��nQ]̈́!�������.fA�@� .~�}�k+����s�:�~ �pW����H,?��eV�0l���T�:\.���"��7#��Y��un�/�k��?���R� l.2$�3Z�Rh�^�@66�h�����X�����D���O#�����D1� ��.��n/R�96���I/=����9�eB��Ci�i��R�]p$C_�����j�\����e���R�^>ߖ'���s�F�'h|	��s���=�/� Y]U~q�HͺԄbI[�=0�w��uf�@)I&$]����+7�(	ʇ��8��ĉ�NȒ!�p���2>נ���Ql���9�芘?�5J�`���I�(�LX9������懻ށo���p�%�������f��6���@���[�Ps�c�"�9�n��y�T���>,�8��=�x?��A,d|��E.���^���*=z�I*�ѿ����g�U㙈MIW"c~C�u��W�Hf�$�9�`���o�!�f9X~��S4�:��pJr܇;�>YR	���	H�#w��*�:�EiG��E��Pw���P��x��7�`ޙ�̔�Je����I@�b�BC���@�CCh�������������q�Z�a���Vc��ӵf����;+��v����{���h���'���Ջ�ي��G�LV.A>t_��u`���1���xa�-���*��|����t`}�7��-\A�N���7�#T���Jjd�O�/p����F�bW�9$x�[�낙��N���P�ao�Ę��ぴ!N���
dպj]�	7w���1	ۚ"G%�c��m�l�IcOo�W)���y��R<�|�������sodZ�4�m�&6u3Wg�dp!�[�;%_Ւ�8R���m1G񔣽�`�(ǖv�$��b��`k{۾�U�CCeY��8F�sXp	�0Q�)�\/�*�.`E#3@�?��d	��*(xH�>��٫MB��\=
�B����i�+��-<�H�ӻ)|�NB4������[^��eH �L�J.�SpO�����냟t-�
�:_BM�0��{�Y�r}���< �E��m����<�A��v�}��U|��ͅ�O3����1�5s\�?�^��G�U�vK"����/��?����Y	��% %�"�9�;$�z
�_�W%՛�@�6�5�ڊ4I؜�/�	�&�*�3-:B�K
�)Fl�;.~/싧p�X��2���Q�W�V�~N�m,�QB�9��aJ�Z� �!F3�[��)��8��?2��Ε{�~��J�W����߳�''�g"���8T��~_w��~^מ�U�ѡ%�#��[�˷d��'���F:����M"�[�ϼZa�ƪ�/3��(�PZ��Ǐl�r��&�u�d4Vf�����׼T���`J�B�^��|"zJ	_�v�!����X�+�h���Lx��p�kg܍�=s��t�C^U��Ȋ3�b@[�㩙�|wOho�L��
a�5I�Oer���E��Bu�E�\~<�=��|?/��DnO;��A;~c���z�ߨ/�"1A0�JY�hRrֈF���(���<-�rz�XP�:q`�0�[0�z1�s�OQ��}��8�`�݂߁m�e����Q�S����Ɯ��ʳ�/M׃6�`{������K���Ýi�(�Ѱ�|�^����E~���YA�X�i-�_�Q}G��x�����}�������0�v��s��1���p�ȓ+��,�Y�e0*]��y��}����lzuؿ�1c�ݿƦ8e�b��<=�Qz,uP4��X�kB���`_ҵ�սC�U���6��%?
օe�9�B��19x��	&۳����x-�v�f��Gnd������I��I��u�� �9"���)�?���?��`�b��TS��0�R���ڧ����u�ŉ�ƃU��O�V=i�YX%�pg���²�_"9���o��a�\kl�mo���4��>�4dO6e�~�Ͼ�F�r�X�Z0������/��[YFޔ�ɨ��֞�	?�V��ާ�X=sdo��_�v����;kt�>_ks3���4g�˘jqWD�,j���RA(`|���ӏ���K��s2{#����
8�
�=$F�jT�>�;���W_-	�*�R����/��/���6z�E����z�:�
��}/��1���s�A��3v��n{�ͻ�NJ�l\�Ԯs����U�'�H�^?�����y3�`LK\�����̳$.`��f����0�n�6�e��ᾩ+�G�_�19¹��`�zdQ<!����Q	�-I�	6ݴPy�i �o����"X�!�{��Z%p����&�dv�)�5wWy
Ѷ� �2l����E?����7�0�-�((Z��-��JڪG��LNo�����������Zn|5���$��,�U(�B�K}���&��d}�+l@<\7T��3E�6���I�m�<�Ć�m�%�S��ar_�;}
a���P�ŗ����ɔ�	��.��|1��f�I��}�H�i�Zק����|�ʛ�L7�y�t%k��vY,hw�K�9q9Ĳ��Y&�h	h����Ё��5�Rp��,ͷ�ڡPӫ��稐DH/:��w$���/�����#��1��k¦�`��rk��F�)���b�&�C9�Y�l���%HT���z���My��-P,s��R�2c����!���b��Q�m&�{� �@��DS�,��7.��G�hu&f�G�&9���ͮ'H�$�R;�_FE��	�Oi�E=7��MG�Ɓ������CK?���0>
E����gO��t��dޟ{H�/�jcJ�sr�!�Qr)M�z~+��A����7���l�,���0�|rT��2$ށ�]E�B�.}Zܒ^]����<m8�5�7� ��5ťL)��
�!�U}tR��G1�ѳ��O�H�����߾/^���7���ɗ����e�`q��;�b��C萦ik�)�W��C��#eeӼaf��Sx��������3WJ��i�*��n`�}�����<�k�4`�xŁ�.[Cv^O�¤��47��1,w��@�DTO�r�zp�M���W�%WX%�;�f��DKn��P�>T�/V;�0yg.ݥ��ye�z3 �7$�6 @�x��a������#C�����@�,��4S�ԥ!Ê6�� g@xã�w����K#GjY9S��Hԗg��M��R�@��'�
���?H�*�t�M�b}˻�g�(����c���l��:!G%;MNr_�.�����Dk���V�@���4��5�M��Pl?�Nm�3]I���H�`_{�1��]F�	(��u� dh��O��#�\c�
dQXVI"P�@��.@��o��N�5A��..1�9΂��O�l�-�Ys8��Rj<��mYKtHi^&+$���/݈���"y6�z���UJ�ʳ��3A�\s̏�"��fE�lh�x��K#�uK6���|qh!`�}/Ė�j��
X}ɽ��׆�4GH�Rq�
�/2~�ˁNS�i����|�É�K����4v�l B�W���BS����W|�%=ӯ���kR?��]�8c������R֜z�<��ҵXoC��m���ŝ;�-Ȥ�[�"�M�eQ��:�J�/{��Vz\2���v@�t�9�"Ђf���㵒���2:S��|--v��1�-z�Ζ8���2��M�}�R'Q�uQ������jv-����%Do��]5��4��s
�B(�I�z�����`���L]�Cy�Jֳ'��B�%EE��e��1}Ҧ�ļ^p��ҍw�Pӎ|�m,+�kw�Nd{ez`ŗ=��0�!���j�w���4B8����Ԡ.�I�_���e.��mU�&}�X#%�i�r�ps~�<m��o��< I},پ�!�쀝����
�^h8)Q�s��bP<��6
��}~
 �fyyxQ0n�\"��ܴ��F�xa6���D�:�i�	+�Te9���@=�L��65JO�N��nf���_�W�$Q6�(5E���=��Y�\Aҡ=��&�8�p����)�:����p`Be�}u�bXT�r
��J:�"����P���k�?�	�+�7N����j��$.���ju���Qt��,�s�"r�
R�7J��Pl��s�ʣ8;��� ����W�Dl<�?b���y��h��gȅ��׆�
��δjR�:AA=Sx�$=n�Q���~}n.�|��X��;>�Ȥ22n��A�r�[�o�kU*�L)6���\RY�J8(.�B�c��j�[�O4�/���}�nk/��Sy�J�Ə�������ҹ���&o����Rj>�ܔam[1[_e�끕��m�J�����/˹�}c@�o���¥3�+�p�J�ifWx���<���@�ɺn�Zp���е��Yo� ����rHLn.�ZL���^>���y�ٯ>�����W`�:	�s�3d�]���OЭnޱw,���Lu�IM�����5���+�>��}12#.�#T}���2.tT��q��`��o�4��᝺����Fk��l����+�����x暔z(���O+����f����O%��%x3�X�_�}�:9�H B!L��=.����#�2o<�lbx�����j��+|�# l|�p���J����+���/�U{O�`�2�t83���iLM��j��M��ԋ������+ 9o���hULGY��ݏ�Y]1�(5ar+�j)����6f�#�)^W_��=b�0t^L+�t\�:��� Kbcm�&�RE)Ƕ�c��_B�v%9�|,W Y3,_+��M=��
��a��#�Ls�9��6�M���6X�=3����#k��;��`�+3�6_�.X����Ԩ�O��U酸������l��?�EP��83I�~LD"��姭2��4�v�)�͞ͱ�={ސ�,�!��6X�	�k~u��,| =k�8IU��ϼ����;���f}S��'�V�0:��.���Xe���;��.9���o�8��K����|5�X]F�pn�i��Z��ɼ�)P�Pųo�6���>67B���p�у��k@��m,֗B( �#�;�]��j�Ր|7���<yK�b����g��~��5$���q�z���J	I����`C�n������Y5�WB-�9F�������ܩyl�Z�)	��M�9u��o�ܔ�{�ժ��N޽���`��i���}!ɫ����@��D
젳�Ȍ�m�:5S�X�D�ڒ���4Tb�|b.��Of�Y�l��bJֲ��W�2)��s~��
b�2pAę�wR���s}ՎT�-��%�F�Ys,�"̊�t��'��E*@�>m�-D�/�ɵ��E����f&N��8�>WJT�P�	�w�4�`C:��vA��pN�[7! ��+6-�Eo�m��`��Pا
�{��D��L��E��Uy$�����}Tc�Y3�� �X	}�mq����Imv,���+�h� ��6&+^����$<
H6���k��(D��^�j�Sc�,�� �)��Zz��hnd��fpo���Ѹ�/��m���t9�M�kuF������׈[=!v%QC�pp}���͆�(�������� G�sFb<r��wPK�$��>��u�����9�PC�y)!B��A�	@�"sL+�s��[UW�?9#oG=}�\��E+l4X����\9O��55��X��,�����s/�����G`�܏ujS�Y�7S�jV27f��}����
�5:�SD	��t��fѼ��N�_���l��D�3�5?]x_��u�O�ȕ��B��u���w�x=� ��o�
v!����]�b�T��N��y��}!�[�؞�l�]Bn� ��gFjr@�b2h��B�Ɵ�m=�u�����զ2CFv�H�7�7�]��A��B�M���fAΛNɔ��<�BEOH�R�&�E����
q���u�M�w���}�C9zR�F����B<r8n:�IQN�#uf�t�Z�$S�m�#�	>=خ���O���ϗ����=)�#+�$Y�Z��͇�c�2�O�R��g$k�j��޹�BP�t��< ��]� A�Ÿ؋�߲]��T��<j��J
4�;���V��(*���&�.�<3|m�[!�*C8��	!�/�$����Ȋ�%F4?h�d�Cc�24t7dD�Z��
��M�+ν��w��v�`���B���b:z0a�ݾ�M�|(2 \50��´�g�4uzTvZJ=�r�醻�]��;�c"�zd���bR�K����8d}�ּ�DEdo>���_�$Kk�C�y�P��{����cɷbr�>]%�9�'�Ѫ���MX|�__��i���8 R6�~P]^�t�;!.la��}j��z�95�o{`X����؃J�9:2����n�ݓ����Fd^�<���~��X
Eb��� 6?O��<��LP-�̮�/蜱�	�ll�v������vv�D�:c|!^	Җ�mݞ�:�:= �,�{�h���'�)�PO����}98cFf�*a!���H�Fݣ�Vܫ���9nd����37e��JSk�5��g#w�������c�z�qZeM�O��$��n)į_,>%�x��W�x�,�QA݀�#�C�ZB��J��� 2�ai�ψ�|��]�$g�+�*��[�nxœk�o�b8�h�zK�ݐW���	�x�pӇ�q�0�޽��G�������ȫx��x��t%p��Y�I�J���-R�o�S�5��	D|$��[	z34J7[V��*U1�l�,���T�D���[WElhLOɪ~���nG��5u�{�Mm�V�F��`T�zFp��4��_d%��C�,��TAdv����Z�kz�W�/�J�	Xz�=�v��2ْ��2�i)C��'���VBK�^2����NZ�7��J��W����w��C�F�Dɳ_��*�W/�0~�uu<��k��~u~����
;6�8�F3��[I�1�ޓW���VH;3��,�z1=����O��{���/W%L�!k�W�[��&�[� 5��L�l҉���4���4X�d�PЗ�c���?,F���?��C^N��&/]~)���������H;��n#XYx�܆0'�D�S�A2C	^�H��M��IsNx�R���\�km���o������aXA��w֋QA�Z�hM�C8 ���<_ ��;r�!�1y�V!j|?��-��x�o)H9[��aI-���2��!��\%!������N6˼�2�z�� Hh_�4�۱(��WS|3*�;}+������ut�Z�_�a�R� �����_ܴorL�D�`�[5�`[�;Ԩ(�W�UNuh�\0\�g��o�P��#�辐B� MȬ�f�i<���`�. ��. �n�����+b����i�I���C5��Y{<�$):�*�	��N���x�_���@�-eD�S݅3��~c�����_�,J�.��R��$��ƲT���y2��M��̱#�ˎ��������q����uD�N�����O�^5ݣf�t$&������T刵ʞ�+^�z�t���*;;��J�b��b
P@~=��o��9$&�o��'�����5���;ޘ�:	Y;��Ei��G=�fy*q
��K'�+ߝ��%J@Va�U\胈r��-��N���h��d�yZ��7�C��!��I�D���݀�+-���.�Ȏ�c*�zU����Q�5��ja%k��Z�]���c��2e݅rU����/'8�a��<W\�)y���io���&�m�T�6 MT������e��K~�m��-�. �U,n�N�Ҩ��Qx�v��N�s
��7=o�TI���<R�!݀�z�Dt�&�YDP@� ̨��1��������*)d��c�� ���#K*���ѭ�D��:Sw�Y9D{o�.]�Q����VP6�6��
~�k�|��Y�j�̋�1q������� K���T
$�4���`������h-?��ݻ��_��m�z�fg`�As�~'L}7���ĶKQ�c*m2_�y�9km�.�/?;�.��~���l����U(�㯋&�=F��e?��} �m��W w�%�pX����0,�����T@�^���?:Y�eRI�9	����sU�ᪿ��'�_��'"Z��M[ǡ`�[t�Ī�Ĵ��e^@m�.ek$�?E�C�fP����ֶZz�3�l��gf,�����m0�qW�� rL,����' �j�:���̢�V����ȁ�j٠@�Ƕ�������k����,�5+n����k�YLv��儈��L�;Or��1w��i)�^���
�������K3~C��+�B� הomD�:A���[j�s���Ϲy��v�N��<�`x�Q�Ϗ��!rV�Kٚ榪,0�n�����@&�?&�L��5���	�����+��sp�Xw"[dx��q�+u&�Ȱ�@Қ�Y��[V?��}� K������k�A����9ͺc&|*����jT%���&.��d�_+��'Ң���0�,��q�������w)�>J��"v��S����"��45����C�Q�ǹc{�A*���Ն�'�q�a@�3~9����I��g�R���ra=s�}���3N���wE�זH�Q|���!��	<��JI�H	W�{������L"�� 
��"�K����z����c9��g���p�%�C��P��8W��:F�������� ��o�^4	egA�ƃ�����s��)L"�R䃕m�1mzaa�XD0\��S�B˥Kk��iA*��w�mZ�L6J����f��G���/��_ȓ�]���>��� �%�;��T}���i�N�I_>h1s��Ԣ$��V~�Hf�I�t�7=�z�o������+�V���1���RztM!�e�Ύ���J��D��X���k��	�/>��VS���3�V끈��fsvxy|�1w�r�*Y��(9?�Ε�.fFn�\}��k
э,�r���x��o݋0�@iC�e3Bx�Rc�o��T�6I�ʍ\�ƖW�-$6�@��1���{�T=H��eK�X1�c���L<���{�T��vr�.��@?��f#����Q�˭0 x�ڮ����~yRʛ1h���TO��Xp�,�K�`W��EW�|G2٪hFu09���V\�/W�Y0Mv�V@Ur�D���C�ŀN���olR|l* _���� ����<���yP����6g9l�3n�\���inAx�8�/O�{��B�KZ�X$��Q��MD9�ޝ�l���ըǡ
�H�Ķ���(��O������xM۹����)�'3�7�RO;�I䭒�	&@<B�0|��3t�U��k��(*���M4�G���#m�������g��v�p�$j�����DOo�O�~Y��#��F��#R���"Q"�d2��P"�]c�J"��,��x�n1�^+� ��E�և܁����-���rO�<�OE���o�f�O�/�i�P����m�G��͔hk_f{����a��|	��oH��tМ�p~,���k�=o5[ҁO�ᑉ�Ty|���^�����08|�?Au��.4+��Ӧ��zYv����{��G�C��j1zgVK��d��"$�9�<��@���/雗�^߈Ǿ���wx��N��y3`��Rc���J,<PM�O6(�>99��F1{��uT�9ڸ�s�i@,�Җm��YG#�tyb��4g|�[oJ:@ش���;O@�&ѿ���<���KNgF����b��pU
�S@O� �%�"�p�r��l�;Ŕv;���q����%�a��Rf�U���V{��.�C`Ac��χ�܊qi�QJ��Z��_g�z��R�����-��/[�?�;a�q����'ϗO�}t�\�q�Gkp��~��mc?r��L���
Z���_A��@�!��*y�a�ƙ�r�9g��'��F}��)����<\��$��8食�+D�������Z)y� 'WB�N# sJ0�����<���7^�l@��0y8���u-���z �p.��%�8R�ϯX��Z���$c^�a�6��[SWl�8�Ģ��3V�l�����ǆ̃�c��Y\_����(!��Y���
�m�˙����[��q,������ESDb�{�X�I��@̢��'	��ӻ`I!�h�B�׉¹H�wi?Xg�ٙ�_�4���o%���(5}��<mb��Z��ΐu�&VO3Ś��ԋZw��`�ޱ�J8��<߮�^����j�+� ݊����X>�hxF��QW�h��nԷ����\��U��Ɨ
�>p#�{0� Lt:!�qO�����K��@�i���\�C�Of�w��V3�K����PŽSx�n��p��!�v��Ud�%=�(��Y��m��]���++�j�2�l�2�ؾ��Ş5G0З�Y��^_��!c?���7����D"�NV&�Tl6� B�4�q3t�"��l %r�����ϳߣb�ZO�-{�����K^p>��Ts���!_��#[ox����Ψ��"Y�P��E�U�-�ɋP(�n��3���?c��4`%	����Mt��8�������ӧ�H�J�L6uj�q���OG/�P�}�ŗ嗌����������?Vgyc^��ް�y�F���}��4W!��՗��/�<��&w.���M=aC˻0��X�XgЧ};̶�b��ՉP�yOn�HJ������n��� I�gt�a��y��t�:U��L����"Y�Ο�Y/u������9>�v-z��Q�m:����S/��e��)�����>Vv
���9��������|�ǔw�I�S�����2�o ���'C#�c�T�5_���0x�߱�����{��B�x��k}x��5��W_���.�y(	.�XRv��4����n�(�E3h2���L�MT{���Z?��^.�qh��c����èO~��N��x��J��(����6?~��U/�µE�AN�L����c~�'�ΰ�b��T
5��y�I�4Ei��pJ�[��EOG�n�����l�]�������tQә�|U��?�9��|fn�Ggp/x�P��73fY�T9X~&DȨ$��U	^�M�5Ҵe�eY�$Z_g�4��x�ȪU�`�D_���)�{�r��n��=��{F|�u99A���YW�B�g�tO�>��	vak Rv�G&�{Df�	�rY�ku\���l�Yu�X�>���ׅ�P�4��P���Pkg���g7=��5H]�nc�xD7�~d�Bb�����XE�E����+ul��D�M^W�B"f)��*V���UmZyv�\��m��>���]*	��_`�ږ���#Y��t���e�3�v�/�#F�ۖ��!S~M�n����#|��|�pL�_��1��dƏ:h{6%ڝI@�{����(�����A�z��� ��݆LU�����_��E�{d����lZV���]�ͤoގ�fX�uL�e�!��H#�3�yn�ӉI�w"A��������:���T��1q�A�`ϒ�2e�p� �q؝#��ØڨD�pfr���j�⎏��hn#�]������{�y* +!Q�026D��A� �k^42Q]�"��5o5�Q����U�CB-v��v ��sYg�V�͗A����4�ڭ�tR3�Oƹ�a�?oF��(<uZm}��j⪚X�!�@o�C�H|+I<�
����G�����.���M4G���`�%��2{�<2����u���E߄%r���IY�k��Y��=������e��m��Va�]�>�L���kIm	�Z��܌��IMl�7!8)gE�tbدJ
>�d~�-J��h��s�ߣK�.�X�+��� W*�&�jH5��Ƚq�(��ǋw�{x����^7��y�1�.�3�ֵԙd���g�U�q-aiP���1� �C���X+��K	cL��:��&\F'��O&$_�ƥn��O��X�H��w�@l	��ro�G��o|DV�S.\BMX��惛ҙ�_5��
���K��غ������c�ݐ���`Mf����#�K�z\�����ᤵzB
/���$�~|����Op�'�ɓ�Hsا[�G��wE��;{(��a�'��zd�~�'0�ܮL�1��^\hjQ	���FyB�,�'e����K�=�vu��+-A�#J{A>:A����ХX�����j�^�?�p��R�B�^�֍¦�c���%u��c��	�!e	K5���˙����:��� E 2m�h0�(٤�n���2A�!a�-!
�i�l^�Q|_@�_�e�L��E�Ȑ=�������v�i F�S�r�Z��q�yp�2Lv>e�]59{�3��������͵�{��r�Dm���tyV/�r��g�TY�ؾ��昕��"�0u�l��_.����A6�zR^�5����!�Ð%�Yj`�jnmS��Z֩� ���1͜����Z���0�N�m�1D�Q���D�L3#7Zy�`jZ��w�K�6�Y���_�#=b�/Ί�G�t�'iĠ�V���-��8��+]�d}��s=�8x�5��@x�:q��oRP������-2T�^�25F}:P���_d�l�9�z`}�Ӭ���qnC���ز>�����q�3�;)+ُ�٩��UcM��;�ܫ��0xy	OY�W�H�q���h.a��� �\z�Β����ot���9�͖�.�۴���<?Rq���O8ڇ�E��Թp�:��L�:�x=�{(�����ҧ<(����/;۬�if�	=�(`�*3�,J^������4�pA�]VH��x���b^C�"xX@L�)�ل��qF%�.���K�����ޑ�ʦ]�m<�sI}X��$�E]S��!�.��U�r=(�5!�W��þm�M2p�;���:�g�<5��R��/�8�[�ݪP�>����}[��t�{��u����kV,3Kb�%�<�Չ-	2�����mf�@��͔�jʈ�:�o��?�K�#	�!������V8�̀������Θ�}�1hڎo�Ɂ�D�a#�<-<6�2b.O��U"RPr����l��(ͥ��>��uAe���I��	�1H��r��*f/��,��8�^�����Hk�)D�=wBI�5ɛ$�:���FSn9��t,�����	�x(�d��RA�􀮈����li�-ٖW�ޅW�Og�2%�5=��8��	�$c��{�@�U[vZE빋���HC ���P{	3��ڹ���W���=���z�c�{%9��3u�AV�.���db��7q�q>�	��E1���|��aF�9�-)W�8;u"1P��ܷ� y	C*e�\�
]���؜�����eH��5Jպ�	�B��#B/�J>���c���D�x�X���`v�b��cŪ�8Gױ�J}���_C�~�,6S�����zT��fӶ�Qv�>&�k*���=�\s�l~c�R>7��P�	�vX��(s򑡼���H�ńwf���}}����w*=��6���F{�S*۲��;���nB��W�vH�teۉO����/#D�ę����ĩ ���x���T(�)��m| 8o�@N�H����QH�#��8�������u���n;#��h�m#ʵ�Q����Ɵb�1��-�a꫼[z'45��׊ ���L�H~c��@Et�Z��%5��6���h��KR�����j�;XF�S��`>�jjM��_���a-c�ц
M�ïxl�:���~��;99[t�Ji=���]4��N��$��o�j%DN��$@e��:u�NK#~��^��z'&��E3�; �`KB�Rr&�����YhԤ���F4L ��'��FU��~�%_Π���4N�΃���=�P9L���������z��6����jkׄ�΍��z��x�0NKœ��O��A;İz޴oU�Tz?Ba��͎y�dtj͝5zX�Fa�u��H]��0�_Z]%̑6�Gkz{�h'���%��FPMJ	v�0s5���j}Lt�kE�yZ��\\�;,�-�S`�\r�drv�q�W;+栧$ߚ,����� ���������WiG�x�A�<	84�kBDe��OBo�0�o,}���?���Ù���m|ZHe4����)f%�i|�r!�ڸ�|Lj l�J�}���q�%���C���e��
E�����Ն'	�܉��}`��j
ЉWEz8�@��}$�	
k����"��q�����V����6풎CǤ�u�����aN/2c(v�'��)��
�˺:Yh{�$9�Hc�&�~��yԷ.�	?�IȒ�{��Ms�}<��	�m)�=�E�93P�LJ�.'�V!D'-?+D��� �����gc��|�`n(ڼ��8A��GB�7�����I�e��$�\3��P��;#I�_SV���"��"gM~ N�oٔ����[�'f�_�8�% �[��u�d6W���tlw��A,�jG���.hȽ���4����w�W�ۋ�Ŧu��X��e��Ѽ�?�O�F S������f-З���[ݯ�ecր�*�n��}[>���Z���K���ƾ�CC��,�E�s嬠ʦ�\��؆O=�P�NV*(Y�9��Z�D{@��x-O8w�B\X�q�)��}Hz���h������[nܲ�e����rIZ�qyF�x�~:��Q����<Y�+��.t P�O�=�A��	�K��1ѓ]C��C��Lh}N!�Vx?�dPޏ�.]D�����~�E5��Oi�r<��L,��w�3� ����\mB1�V���F��ڰĊ�AR��dY��}�F�E��o6��2`�z��E�|η��w}1G<��Y,�e�+���+#�J�7�?�?�͙���27X��WN��tz�( �a�������r��~�J���QMT,����gw� ��`$#am���li#Βs�D߾�}!��"�L�>.�!E����[�?#��=�d��#R� ��;qO�������f�_���Y�Wأˑ�GQe���\�k��m)������nG>�I>��x��1�������)w�[b]5���c�UYʯ<d�"��yDF��$#75Щ�b4�{�R
�&\��1$(��`Fx:(C�*�̝�I��\���7f�F��K<	�#��j�BeۈbM|�x��?��J�̻�>�?Z��E���j�G}�ȵ��bC��t s�$L'����G�S��UC���N
�=z�>	�{n����K��u	I>U����~!L�kr��s�����Vj�~�[>vS&�qNxf�U7�_�F��TгN���0�rp��H��f�1
�g��i{������A�әb���n
1�*��S��h�-�_�Ƙ���WB����UH�p��mL�\�
�{o=c���d���̦vI��H�v�鯨Y��ap�j�
7��f���m#��9�� �Ɂ\�1#���ۿ��A��$��e5���J�"��R��S����[0�)����:�����'mF/1��A��|��~��7�P�6Z��L��fy~5?��d�����5��ߏ�D��r䀽e�~-�ƅ���D;���qd$^p�b���~��BK���������6���F@�����ʓ���Rk��t���N*f�(���u0�vl����D�=��y%��O Y^�����Ъp��~Ɋ�J�������y�.k��Q4E��'.��&ʽK�
�f�Y����~�e�Ժ~Z&�N���s�����q�"C��M�(Q��Cwױ�q<T}A���zG��X�ř;�-�t�{} J�·���ƨ+�n.&	�X���Y-�ǹ:V
r`�R�؝V�]�ݷ�k�1�z� ��ղ-Ks�u�2��_���ݾTT�ܟ�)G���\h� ��K���YW�4�/�����ܬQ�]�S�M
�[��G���.R��6�_��!v�m�u��Uj{�@���7b��y,�� t,�pM�2ќ��Ҙ��.�̔|S�Wx����R�p_s4Z���>;E�����e/V�5q�#'n��#6k䪍
�n�$�����i]�0�O�l%~�^d.�J���}��H���Mk�c����w�6G��ߊS��Ug��6��&�����{Xz�M�l��>\�c{��u�,��i�yL���"1,NeK��Jλ�"�ޮ����^h�=����*O����,rY>�ަ{.��|6z��y�H�d��3��IĮ' <�?��0����6���g�w��ROxkF*@��0�[՝�=v��ɹـ�� ���0���M��z�=�v�_�>}ɫ��AɯcͿ�M9��Pc4@�U�﬒�I�IF,���v"���-�N�e)��"����E��ؘV '5�^��-�q���.���#��s��1�E�S��-�
yz��)�ț�X)+a�[��EG�t$���=��,	{��u<d#v�s{��yy����`��T=c�}m��D��K	�I���xϘ�ج�� H��鐛(.�`�vT������d���!�����8�*]~�����^���w̮)�^P�������〇� ��[~k j�E�z�#߉�� �_GZ��)Z4!@9�����3!(a.�z�#�����[ˋӄ	�8I��'��L�a��Bu����l�?��Q�$J�U�������k!�m*�ϗ�yN|�H(�ǰ#�~��V�bg�)��u�F�p�kR�J�3����1��u�	6���E�%0)�h�	�����<&JFQ^'xuO%�C/�3
ǯ��������I��#X���!�$ӛ�VG܈"v��M�� z�n܈8P��
�Bo�t��ɭ& �L��u<A0��V��o&�N��ެ7�G�R) i�Y�.{ݺ՟�-�m=�Hg\X��F��ɭ���W���蔚pLd�1l��s��K�kx�,��r�����6��K>���ݼs��y�J�M�L�k]6��V�(��m��(� 
5���&��5�6i^w:<w��1��;��&0)Le��'�={#�܄ bO�qTLP�u&�jo�3�{�T��������wG\)^+� ���j����� ��}�i^|z
)[������&J]��n��Q���KeD�O�9{A���N*��s���ntH&���E^s�<����aW�n�UlX�	�u�}H!u
l�to܈V�j>Ԥ8� ���eV)m)��R�O�L_�.��`�ҢjV����M
�2�vСR�U)��{��d��]��7�
�)`���Em�@uȖ�͞�V�ze�!gN�,�?�R�p�dl��""Oք8%�JcG;�1��a��r{6�Y�.��U|�f�����4%�}� 2ݾ"��
��-l�����W�����}˃ӷ��׷
_C<߄�^�z�8õ�z��A0�:�����������%d���}T@�>e��mz�l9 ���vA
�of�U���A����ܥ��y9%�%Hs.9rV�bh(��_�4,iF�@�D	�0���L��h�fT�Y#y>D^�1);�N�	yk�a�,�+���	hև!,%`~��ٿ���^�>��.fP�g��e��R����7��G{!/�[�'���]s�׀ׁa��Uّ$��O�Y9{�M亁Q�=UwU�6+pW'�2J�,���=�ް����v���I	�;�矍�1���Ҍ��"�3������~�s�k��G�gl'�Guܰ�mcŝt���.�����k�t���%�M|ѐe�X��
���M"�!����2z�o�������:o&G�0xV�k*��h�1��}�$T�	>�W7��}i�W�?:
��L�M��x��Nj��ԃt/����թc��V��k�zm�da*^أ:ܨ�x�R�t�w��+�3�gR����J���6zc�����N�N�N��N*է��.�2\���Wm�����J��re0dc"�
�Z���蘞u��� 	OvW�JZ��+�G���V �"�S{��C�
�L�W�\T�Ъ��T1���?�Iwjo�`b���2�Lz�����*�r�=�1]g�>�\�*���c��qd'=����L�#{o6���(�0�c�[}�_��鷀	j�z�(���2�O?���L`�6J�u�)�+V��D��ԦsU�������[b�	�ɂ4��m�A]W��?&� A�:c��1�4罨y�kS%��Z�4GJT�����D.0�u�k`�5z�pV��%�1����N�i�荕$��v*��٥Ŵ��ؾ��P[��
�<c��|a�c� �;��CÙ��?���'�	I�o��m�'�p�|��"{Lz�)h+kW8h�j��0�?W�_/��Ǩ���LtZ�l]ݞ�`��n��2��+�*�{���i��r*����H�w�6"*���Ź@��`è��)%�ПaW��#:}#tQ�7��V� ����t��d'H��G�e��.�boK	�i�m��v��[�T�4�~���U�P�K�U��V�X] �h��f0����x��?�ܩo�s�'�ۣ2��"a�K}ᥓ�p��-�N:;�b���Y	�+|K�zt����[g����t�RT�zj٢Y���`�0�jh[J��2,�t�h�WR) ��0(z��m�5�xuƘ�_�>	�rNB��0���p����.wĶ���GD��s__v�K�:��[�1l��.����4�T��}d��?��(�	����OlOȳ怔t���GjV�LM䶱��O$�ݳ��W��vl���, �Y!�:�&�THɍe�p�By��G;��)�0�t��������8�?�D�&t������#��\�M�������/���a�FLA"�B��O��gМ5����t�Yx�;�Mq�i�[s+�_
H��I�[��WJ� ����g�F�+�.��k��6=�b&��͞T�S8=��B��T~S�|�Bn��3}:5��f�s�w�d�@�u&�Lg��
��Hb�7N@O����.���/&�,���� ��1n�Hԋ�in���4�]���C����`�(��Rmh�Fk}&��M��#Ո��c��*񢿣�T�9߿�����V���g؝��t&	|Ԏ�r�w8R_�7�R�rU���wfQ��uG��=]�B3�7�Ŝ�#��Ŝ��1��LMI�Ȑ/��C��D���W��ǰ��x�+q�6�ӟ��	��G$�#�����!�����ɬª�Y����e��% �2���78w�����Lt���*�
�zC�,�Ԅٯ������Ͷ(��z8�~��Ro��)�����C�^�ɤJ�������i�9���jnν}�6bi���[KGMB)�LcgxGܰ��u(TfH�8B���O���tC�'-i|���$��.�֣f�V�����6~���'�f�a���h
�:0"�9�9���R���P,�[
�|'��	�3-Т�7j"�D�4�4FZ���O��O)e����/��ĸv�n�!�Cm�h�Q�[x�����ѧ�(x_��Y�"�
Ԓ���E��=�]5%@����T^�qsA 	_'=����Ӹ@_�f�fkz6���j��@���선���	�'����zn� a7&��O'Iּb�L�۠+���ց��#+�Y�[lJ�����	��G2Jt-d���.9#�I$�"5�c�Df%��d��9T�K����=~�˄�h���o�e^�?�}��7�_KR�I ��ր�r���}���"�l����x:������38�I�����y"�D�{���/��Qß�J��$��֏��A�31���O����m�q,�����2h
f�l��'}F��8M��t�v+gϼ=^�)Q	)�^`�g����SDcu��BD[��CYͽf(���2�j8EL"���)0��xM�5�c�f���_a��ƧY}���k��G��Z�y�k�VYz�І�� ��S�c�gX��F秥+�NSc0��Y�~4L��y�%��Sr��ܨ�;H���f�N@��@���{�3�%�#���wf�,��3qa��#kH���o�����/YGIO�Giя`�Xr07?�r�6uH���!P��/��|b�U3����+�>��+`0��wkh��Ws��:�,�j�6��*�v��=7�ҿ@�vO�FQd������5��bĺ�@�]�G�P�{gF��b=$>�8#�G#�m��@���A}��8�.��4YS]���a�{Q+H3�e����=ξIP�{�|�`���*�"q
�@,0�8��.*��	�0	�{�E9�U��w���x�!Ƽ�A��r�B������ V�-�P"Y,�m�֙X"&�g"t��2K�2��n�P(n�ݏ��AY>��qX�)gd�Ki�(^8� �L����JyG
C&D��	���z��u�r/��ۻ���m��WE�r���?V����Dc�<Dk�=_���U{Z	!$VIy`�5$�O�AM�_�r��c]c�7h��`���US
W�NZ���
�m�>�]����+��٠��xE|�"K��Im#����A3�~F)ǝ�(�\��vvE\�-�Eݘ���h�(,	�/H��m$棒P��욆�3��I�i�<��Xp��tu2�K�rŦ,^�~�Ng����+��P�Tɞa���P�XR��,���se�6E+�����3� �>�D2��_�]��X�'B�(�.�SM��+�$�58�5�a`�W>J�J���h����a׆Ǳb����K�����ҹ8'��BBŨS�~��m�E�mdAd����v�zc�&˵	�M�����������63�8X���;�MG�
���M��78�r�*�b���c!BL�|�8���O���xp:�a��P�BPs�{�Ӑv�`��� �{jI�]Ǩ.# P���)!Mp@�K|e�Z_W�d	����f���2��H�Uv��\�`��������q%6ӎN����#yG�
87T	x�Z�= ��wg�pV��wrK��b�����s���{���[�#J���»�V:I�s{��� ��810l�\�e�G�/���'��%���)�4����!�O*KDr-/y��3�h8�:;��\��߅C|��9`��Gd2�" �߆/��i� ZPn��*��F���s�\��J����q�����ST�i�������l/���m�+�s9�8e8Y���=R�Js.�`6j[b#r�v���p(�� ��`a�*C<ڊ-�%R)�����|��F��#��$�i�`�y�ͧ�:��-c�^kVU#����0:������~6��^^�|3�!�
�N�����oWH�H��6�Jǻ;��b�˟�Bm��
A��i����`����O��u7]饰�2�_�q2�L� \gE�Db�r�L�"�y-tڇ�;b@�~�f&�}��Z5]mKL�ْɃK ��ۨ'L�Wd�PS$|N]���,g�4�nA@�L�3y��m �3��*5zB����O�}.!%>vΥK�4�� ���j�6ದ�2���Oܘ��� �#B�(b�$m��H"�d{�?�;\tfͻ릓������:h��2��>��>LM�憏tA��ڈ˓� �Uu��y������ �1s_�dVr���îV3y"i�@��,e���k�������&1I&�r0��]y��>e�Q���_���k��$�=f�s�5?�6C]�vk5�J���.aĭ�g��$a5��J2<YgP��
:�[!����Oz��kN�FB�ƴ����8��j��`��iW΁�M
`�A��/%4�}�t�׿t9���?|f�3�C����}��q�mI�u-R�q��&%gM:+�yH��7��l� V9Ħ �GDOL�ds=<#Q/�z���$/>�p��>�%8ˉ�v`�G��Z3>S��ńOi�9 �֨@r(��o�0�¦��%��=��e@�� ���2�2XG:�v�T�Q�������hi ���A7������5M̡��Q��>F02ꚁ-+Zo�.��4�WM��`lR�W�!|�ۃ穮&���z���H
P��u�s�YN�؈��g|�%��Q<�g�`�����È�3Я�=d���������B�(��oBWɈ��&��E,�%5����;/�+��㎆�7	��fSp �/d^�+s�%�N�U('I��g�P�N�[i�� <d�fȟ�@��G�jSX[�^�{�M���������m�j�"��ߚ﯏�����|���Xs\K��+|D=�6uΦ��U����rݧ1�u���Ǯ��VEP�~`Ο�-�m}+O����Cu�]木���9�#����CM����Zk�&��E�^��7mM?9����Q��Z?�~�5�Z�D	`�>��0���`z����F�KIP����F����s���G����:7-A��jQÕ�ק=^��F���!S�D�`|`�O׍$�m�_|1�~4�/�~��z��7����z�M"������ˉ������<5�e�l�����};��4n�U�`�pO�/@��Ky�X��7f}���/�s	z25Da��/������K��׽F����b��~P�Ze�����ڇ�+�N�w���k"˒�G�M�n�1��9 ��]E�/�	qex�Nu'Y��u{���0o��������O�N#�	��>�}\;�4���9�����L=.�dX����/��U���i�-ƯL���&��y��F�	���k��!w*cԓ��F?1K�SM�l�h�8���0XT��UE���mp�H���W&e�W�$��VS�{�;�TӜ��=阮��.��q���y�+��-C���}%i�T����`欷M����8�q(lrm�,/�+LM~�t�r7Y-Y��0��Ǐ	��q�Vm���+dA/g�:=�����}��S.+��@C�i�)�70��0��#GB4�Ғ;��\쥂�B�̢5)̿���'$N�}�r�7�0�i.���c�3�����6&��pW��Q_&p=̵uq�=N .Lxѓ=��DU�Q�|bC���[�L4�g$v��F,zk�%i��M�A��I��	���MɭM��>�UxbEd�h��荰Ϝ9< �D-���A�R�h��|x�L����@ɘK�6{()�����N���șx�L�H�v���}�"�M�r�@����/G�驫��4K��%
�b����^Q=���$Z��	0'�ק���B\�f�h��!Շ>d9���.�G�F��~�0����yn�I����2%�	����7C���knSۼg	L��!؂θ	O�y*��Xˢ;J�'-�<��7�G�	�y�*�U�YP���[��s\Ƞ��&f����#�
�/�X�k�O�5���%E�����1���!� �:�1���DQ��|��{�4���� �\\�UE�Ai����l�@wĩ��<F�y/��](y@�D�rF�U��#���0G�՘8L�vS�J<d3�a�@B<�=��Dr<�.ng�W��S�J�%�Ra��$@/_�5���xC*-�_tT��~�e�I�8�K���.^�g�d w�v�:��
�a����0��0��f�����c$DZ&�M\t,��e�����:�e+d	�&\2��R�k�d��" ��J6+�u�P$AD�J{�~B�׆�C!V�z�&,=�'�X(�:�8.���Q{���Q>��jj�B��8�b�Cz/'��Fb�n�me��ɝ����Q(�q��f÷�@rȬ��>j~��������>g���]I�a2���)���N��v�6M��%�������hHAY�e����� ��O��Yp���·j�"�|�Y����{��}v�Ǥ����3%���]
�fJ�맣J�ΰ���~x���?P6Z��3I�6~��c��
���R����6ԧ]�w)��Ip0��r]Z�(�uh3T�M��'��q�衱C�f��Uy��P~h�ŝ�!v��܆� `-"/�t�|��|OVR0�B��x_��CO�A�%�j�v!�,�	A?��-6����j�5Y\�ڡRA0͈���v�@�@y��y2Rf�����7/�|Ѯ���d��U��ug�h�8B��qKȣ��Z��Q~��� wWo��}!�)�Z����9�j<~�>諭�H�;LS8h!�OwRU?��/u��2�����F~x� ;D��i���/����|c6s��� � Q�!]�.~�ڇ���A��
�d7:�-P,�������
Ĉ�+�]>����p%a�9�l�=�pۑ<��2�L-���	����ˁ�.�ߌ�s�q\B�P�z�p�����z����뾕j&��@ᴁQ�R���o/�>���ϧK�����wΛM�)skd`����	��:f"cp� ܋he�De�DW�W��
(���M��=J-��uIg�Q�.�YF-����(Y���N)-�����=�j�N����0�8����O|C;�B�dL{�&�#�g��
D�yE2Z�N�KE�Y��B���O�6�e>?[�����`)b^`����B����]Dt�j`x�ا�k��v��/03_�2�)�'� �����n��Q�Ȏ�lځv4|�W��M�����kq�Gִ8	$�H�9�f�u��_���ժu�[�چK����81�Nә�i�k�ՎJ'渐��1 }S�t��?���&��[��p2?&���-4;j�|x`?l~�L����H����9������b���E|
����A2���	���`�8[?�<LN�.*|�������ؓbR�u}�{8�68�#��*~[{�>���� �9(�)�������J']l)F�u��P��fX6�#g��iୀ�h/���,j�w4�Aa�ی��.�JXjn} �s/^`���E�����!�(,i
LaQg��RI޹`;)\�)�������9,��Cﾄx�t� ��Z����m�%���JU}vQ�R�����M��&z4�r�)���H.�"��e\ ��4��e��X�������:���hŧ+�e��(�"����؏tT��y�,��8`=S���g`��h%?J��&cb� ��DGm��6O6 K����N�t�7�G�������'~�h��C���tdz���g�#�#��ZiK7m�/ip���N�r��	G��ڥ�!.�c�qN�`9���c]i����7"�<L�8�S�:$��T!��:��֨1��Q��-����>���zur̯�~��ãK�s�Ts#{#��Q�+�SS�Sm���>��GuXȺ˂Ib��@ 9+#�ЖWf_�����f���ms��nDA���&յ�W��vP�������¨����TՀO�.H�t�C��I��q��(���a�LQ���!3��
�*������u�:���"�%�w��",f&L�-c�u
\K;NV]*��WXG5����;���+�2՜��0˻��M^6Fh$�'J�}񂉿l��w�!R����tVZ'�x�t�"�r��|����v=d�����w%���lo�F��-I3�������1~�`���uL�&��E��w~� �t��ϗ�M+����(��;w��t��_�0���ٙ�6�0�q/��h��$RE�vjc��*�A��􏓇�:Z 6˺2��J��������h���u�|�W�[h^�{��>���Q|�ȫ@��`�|���(�[~h%�G��D�(�[>�B���F��	�;�8h�a��x���4��«T���L�� ��{�㍗�⍓��~�aj1͜H@�`Θg���A���YK����<�!z�������d#;NQ6]*L���TZ����c�L:�����S���+h��Ѱ�a���ԛ�b4=T����UU=�5﬊��������Ot֌)qP��B�:Q֙Yz��A�]@����Ŏ���qs�%tb��ԱG�Mk $77QK���ӰM� M���nt�v{����񢩙�	���-ڱ1���s�ٞ[A���%�K���u}��%�EQ완\x��J��7n�+��<���SI�0a _89��eB��_�飓8y��]P�x��W�
����	Ѡ�Po>\t�\[���P�	�՞'i�|N�7�Ej$x��L�\8���Tr�=Fh�<f:,4��p�7��⍬N^��
w+�Ơ��Os9Nn��8hW���/-�ڣ���l�=� �
׉�_s��1�w{�*Į�Z�G?@����+��eVHX�Dr�ç7�jDj6�(R�c�c@I)����)a��?�FEq����T��Q��ȸnL�c�M}�F���R@�s���!�w�F%Sa�]v�����ڸ}�hMEW�B29��(�����{���;���k;�&��(T�ԋ�L[�b�'>�|f�83�����E���%���
�k{b���Zy\�I�G���|�	���=s=Jy.����
�E�2�%f`ϫ����W����G� e�Wk`a��Vq��,�nF�����8��÷�b�)Hӏ�͢o���8h�}i���(7���W���TH2�E��l1��6�[��/�z�s��}�k4e��88�I�h�D�\�V#��=t��֘y�{��nJCa͟����ٗ!^�=��/��apN�ʋش�R��_J��a�p��V5�1���T{ŐNe!"DI�V����9N�7�u���#{�
�\�cU�2Ⱥ�ٕu�c�b�hkY�,���d�b���H�$o��������f�aA�`�5�1T��ҽ��8$�ɂ����	K(l�S�����y�
6�t.�v��=��Bkn>�}�����{ ��vr��\��P ��xmG�{�	����+
Bt:�j�[yj�xz.f�*�Qhlq�T��}��Z�	�v��,f�r;��^��{�T��{2��Mڰ�4c>��xd�	�g����p����SY��ŐQ�k������\3�V���u��I�.#ψ�ϕ�L��ݗ�*��TJ�iY��X�h�^+D�ɵ��/�ڍ��6P\�.� ��;�(�f��Lz�7��� �Mlo'|���NԠt�����H'�����NK���Hm����QG��y�
��U�Ch�AEJ��8�1'V?�5���/E��2�霰�&����8�%��]Y��/���✛��s�ٌ$1a�]P]Ì�� �/V�U|L���W��NaA�"��Z��'K�e�ȋ{�n�>`?Fh�% �Vb��0������LL�Q�u_|_��kG�O����PKh#��}��V"�)�*����B���X�|F�?g��;���/���g���F�"kQX3��|��Fw��YN�^�Y�m�/�fw�K����Bu��7�~T� �T��q��ᔥ���i8���2���{�
���Ro�Lਗ਼XC�0.<w �����v О���BB���K��*�/���>��h���Z�=r�}-��_�W�7@)(�����
�m�Nt���b$+�!;�������Q�U+�nӸ����������(LC���2[CE�����W��*��ݯ��޴�ci)p{�����	�Vk�c>� ���U(OLgE��KT���|f�JAM ���F"a��A�����k4,�ZL�bYDx�#��G�v3����&�>v\mKHǋ pKgr�
�ˀR�$�j��M�K�iۙ�����,�����8I�Wq����@��	M����@��K�穾�{�x���a�7��a�<Q��q��,2B�C%��҉J�T4�5~��D�]��FYJ��md^k[(�AeV��:�'^%���%ʸ�B,�]�A ��ʖ��U4{-?)�<�d{��*�G#�۫�ȋi�Q(w�($3�[\���e�|��i���NN?��Lj
�tEp`��#D�٫��??7ͤr���s&�V��U'�i}2�T(DHY�&�d�k��B1��G->��j2�p����#M���X�a�����t_�f/%���]fܕ8mb��F���|F��G���=m$�#	tߊ����1Uq�(|ǒ}
PF.�(�����~�_^�%��dKؑh�5��~�G�u����ĥ4�1k��C1�@��%GʕS;��j���*���)K4�yHf����weV�ߨ����'�*1�Z��NNޚ\�B6���KhGܺ��|��Ϲ� U�J�洲��f�m��R=�V�-U�9��t?��[O����"�Z�d�v�I�2�Y�,U�b��rs8��$U~[CƊo� �m�8�����Mswa3��-6�
�7�`�h[����e�͆��{��c?s�&Gc�.�9�$��$Ș��+
� 0��R+6��n,��S�k|86#�Q�e:��[����hD"Ā�YN�B�$���b1&��9'�MBKy�|B:[�I�]�d�U�HqW�8���Rտ�*~S�7�!��ѧJ+.u!�;�n�۶p���p�8�����
+���l���@���x+ �����27u�%�Q��-Hd٨u��=�N%WA�c���?��}G�z�A��9w�ڀX��jוq�)[���=�F�Q�\�X�����j�5芥�P�)�N��+c�+�O*�Q��=��+��9<�w�"���f>�8t�����{yK ��^��`I�9���|g��Bj	�_���q>�c�/�D������@0e|����e�2oFQ�
�oƱB}^��]������e$�����ʠ�|�E:����.%�^�BYO'�Gݯ�I�o	�k��ێ���V��Dl^��i��g������T��7A�#��D����%i�&�ߍȢ!���}�J��#��������틯���D�(��T]:O�=	SB�g?��XCn���/�ϩ������]�rt�/� E�2R,����������rrY���ү��I��&q�Gi�u@���
��^���&'�grq4� ��iB�mV!�~u�iB�ϸGN�@��r�ۗ�-�ۗ��4Y�!up����VX�[¨A�Qa<��.�O���4���t�fs-�����Q��F,oa�3��D�@ڮ(#Ӄ/n����s�%}<��#L��A�P��0�ͼG�x����n�g��G֑=5�ن=�l�z&o�x�45�mm8y0�(*�T�����/8��x�(��'`���'h��mā��ݰ��b؟�O���_���M͵}>�6f�&��4����BJ�Tޗ�h0����?��33%f���c��YRAu��G^ĕs���OǷ�H�/i][E?�z?��� ,T;DC���	�������y��qrk���]�,�M;y�=�!�}YuAe�Eep�����槅��lK
S����;G�L~��?Y�L�xJ��y�R���Rb�3z���ɠ�/�m�^sZ}v�K.{F�б�Sr�s�٦ ԇ�Q�p�s�t��_3Yp��0P)
����jj��=.����%�y�6@�7����Bv�-)�3g��rd~)%s@;��(P51��#ۭH�j2kBs�͖��F�ۍ�~#��U��he�~� �CS:�^9gDѡ���������u�̙@ D/��Jn\۴O'�øI���*z�zs��>4E��h�iP=7"�����HQgW��@��XJ��Y��o/cv�).y��<}���q�j!i0]{2�_vi�:�i�e�NI�M�T�����-	�E��z:��,�����#�*�9�B!�PF�W�����S�F�`>��I���� �IҢ\�+��ƣ$y��R:��z�r��*Yw��!�U9��|Xg_�����S����G+�1��d�2��L+��o���%��{����1���ML�[$4P�e�i��Ys��A�<:�+Y�z[��f�٣%�*ˠΖ����܄V��'��� ��H&�pY8~_�4 Й�L�F�	5h��A�PT�-u�Ĺo-�U�[sk��j�#���`�p	}�*�̬ᘇ'0�����M��0A�bNC���^��;�S�	��r�똫����	h��+���V�H�0U���@;�W�%��7X�����3jxȠ�v�7V]����u��� 0e���u�g�h���C���Z��D�h��>a�w��c��d�����$ʾ�)<�Rm��)'-��������$HV���	S���p���|�ʢp�Dvl	����K�;�IJf`�3\F\/Ue��7	���M����EW�,��T#��	PΒ7��q��j�ZC 	U��KC©f
&m���'�_�=�_�O"ٽ���[�C1I�5�w��#R��|�2�Z��fK��P<r-��o�j��kĉ/�@4�������G.�Q4C/�c�	�p��[i?Q�)�HOؙܝ��[�r����
͕�7�
^�zJf �V�4Ķ��OWV�X�E\���l;-�%0ć�GQ�������Tzj\O^S��#j���Ы�MP7��E���Lj���c��V�c:�
�p��� �;�V��8h,�(�M߸�j��YK�+%�6����`�1�nv��Q?�Ԯ�n�}�]�J�r���c��OTLj_S۬W��'�j{.��K|'�9�,�դ#�&����,�jV�\=�tfF�m��_�s���A��tٻ���w&[37k Pק�b�n�[CY��c �c�p�c�:��gt!��R�ܯЙ@^�,�a�k��\�z^T���`��+��G��N3�}�o���ISD�������Xɷ�}v��0��@���/��JQ��}m�R
�_�}W2�|1������~@ѝ�:J�1W�*���'�k@P;�X�x��-`�ޑI`�����+J�t\��h�Weֵ�^��.��O1�
Y7��`G_>���p��%��I�	��!D� p2�/j9�R:E *z+���*!�Ј5O���+d���=HY7o�����JV|"�Θu���qg�(.�̟����K���� x*@���j���(Ġ=2�D�a�Q�����*ȼ��X\�����=��x�hp܍����I(���@���1�p���03��J�B(ڡP~�(��������-���Ǎ"f��j�)2گb��I��"'7�(�3U��N��tSA��7&�3!?�,5��}�Jim��SU��f'�k5�2G@�E^�v!/ar:b�,�%��#��e�S�Z��Q���pƈyc�r�*��`z�kDO��U�4���.	�N���� =�*4�����"����U�Mo0̿ur�s"��c	3�7ND���j�Bd������0:G$Xd\!�V�g�-��P��M��j�֜�����N'���X�U�9#G����0�2ѽb;Ʊ�E���@ �/���,�D,p�O1= q�8�&��疷�� ���,)ߓ�ܨ}(Y��}��|����Wx��UJ3��!�kށ�
u�aT����;uluno����*�p���E��TCZׇq�D�R
��j]���zxiRz�@����^�Q-����îL�����w2R��jg����"1ݨ���ɃE��S�ƈbay^/˫C)��86:[7�j�W]���_�� ��5Őz>����Zd�X�hbj6�p����ڼ�����h�V6dн�;$u�{��S��������A�7�$^k���h�갫^w�w�&��[�s���eGj�S�乜��,��ŖY>$������,��%��������0+��\��C���EP����z7�'
[!�mU.��شo�Arwh]�z�m��Ģ�O��z�ڛѨ���^>(���,Yu��J�̡�l��}g*Si|�V�V����5�[ꗡN�����	�Ʊj�s��Kڏc�<]& ���f8�td��X�K��:܍_d��A0$�,��'I�Et�P��1�䤷�$!��0�� I�-4�� �.�o�C'>Yȋ���ݱ	6cV�^`���?�m'��_��Y ���Yt��^<=�o�3P�?��؏v��'��ꆀP]h�$D��z�,Jr�n����xu[�QRO`��=U��w�^e�o���
?:t}m{C���U����)-������͢�5L{:�e�������sCF�lͮ�4�� ��c��ht̒Bi+?��F�̻�p�3�W�!�`9t��g���'/��E.TI�ǭ�E�kk8��N��E�\�Q���HIc\VL���?Ѥ���E�Z#��}�"���Ҙ4B$��`���R���!�?�S�ȃ��_DL�B��}��كiJ�E>����	}=`���HR��j@51������k	�~��9�e3���:v� �)��J���s[@o�����q��y�ӐvT���r�@�=<D�a��ǫ�}h"�	�}�?��;bs�P�'�����9U��c��m�\%����U�7�p���#��:/�i�u�Pm� N8�D/`ꅳ.,Һ?�mG�Df9���廖&�nͥWm��jeG�Ul��ߏ[f��ב��%�0�{Jk��L6�/ꍭ҂	-�p�Ok��'UT����d��c�RM��WT�1�{�m�aD����t~� }>��8�hų�^=��q���G�Xk41W��Դ_��s"�C0��3��B)��>�>\wi6G3�Q�����ӆ�zj�,6�E��}�!����ń�]ㅛ��P?w'GU+wU�$+n?�M�Ɔ]�O�ed����V$�hk��s�t")�M�ʖ>��,��Ӊw��d���� ��T�}��S��-tP@J�8@,�4�Ev��z�TD�ͣ|��a1!u][�-lOW�6��R@�������ؐþ�.w+���Ǣ�}j��K�h���;����*�)�$Ko$y���b��P�K9|iMv��@�9椕��M?)�1A7����K8^h$�R�DN�9`ja�����L� ��o?��[]��psdJ1�ڟE �,�o��,@KC�@�"�T�@�-��8����L�.��z��%zzhS v��35i�l���_������RsY���7���+e�)�8�p�����a����c�R+ �{V�Z!�6�󝟘֬�����}P"��M�|E"2s�R�����N��y��Gv�h��W>����toYYS��0>Ma����0�r�/��h���$%���FJV���X�9�.��ƅ�A&�� ݇�U���6&@��U@�]�@�W T^Y�+�v�ʻ��RNJ��I�����39��5�,�����AH3�
N1&
�C�pD����a��uo� �&��o��H���Ṫn�'�����:G�a�/l�C]>Y���&�9̲,�U��. ��,)����@��jxEQ��V�	��w]�� ����ޖ�Tc�|f=�@���e�c�+G&;8y[Q����Z�U�Y����m�X�t�"%}�\��b �a?�j�����������\�y$��� ���rLm������9��a��U
f�_;2����t'ad�}Ӌ(�&�*X����;�_$6����.����$+_S䩐/�f�:�,#B��I���7�ǆ׬ߜ�<t��Q�^��3w쑘�B6�,����~AM7{�H��ϑ;Z���RT�ol���e�8�/iqxt�n.������8��f����ͬ�վ7�I"T� ����ͨ٤�g�1go*9ǅ�q�$�e��ҵ'񾑄�&)ә�I�u��l}��耦�˖��d@��D�,�1��[�2<�:�P`S�l�-�O��c���֨k��@��E�T�x8��܅�o�ذ�뻾A�ף�愤���G	�إ��@����R*M��"S�-�/ٷ���y�}\3bߨ�C@vh�m�{���������B��g���y�6��2� λ�W�%P�6%&���.���>�	{�~4��܃P�%bēO�z�:K���W$�~��}��j^	UKk$��飲b��U�I�~�"� �V'�E�RL�݈v�d^n[�_��U(}#M�uyƻ.�&�<P���0��T!a1���?�u�u%3�D����!3�0T�Vy+P޿G��	���D9D�_��(Fa�.�P���(g��!��T��'"%=B	�n����D��E#� ؙ�

��_H��P��0('����7T�
�(��&C�,Zy�m#zYP�0��޻W,�󡔋�_ih�`�`ώc d����Z��m,!o��!c$���h_a��AD99<Jh|�6%8��zA���cR��v1�|p�����Nt+ɠ�Y�]���	�Zm?��A�|��"KR�����S�=���,�D>H6!�����WM��o�&�v
���v|hd�Tg�ϳ�o��d3�́z ���h�����9`6�8P������'�,D�eY+,����zy�L|��C�
eܞ�Ŕܡbr��>!C���H
~�۪~'���ފz)ؾuC��R#)��*"���� �l2 7<V���6�iP@�y��z���`��@��rËUJ�����P�+��Rnw��0]�J�+0��5��/�k�s�U�߳]�6�밆eK�G��m�Ri��yX�N�
�}η[u����@G�H��hp4���|��t1J\S�b���KWѐ?�Ƒ�g����H��$Qs	T�̳,��e��h��������q������l<֠���_d��7C\���)d62�:�'��w ���/I0l��ҬD�9n##��K�ì�3�Ӣ�6�6�=���K,�5
Ҝ�p��#��)��B���~�^��K�J]/H�O.rNS�F��AD��=�f��@2�T��j�дJ�?��ӀZa��j��*�T�X�V[ez���>ZD��IuF��~��?�+[ϟ|Eaw�Cf6�A�+��/�z�YbaFL��h�R]U�Xߓ7���jX�nh/������LF����|@[�g���+�w����1P%���r3)H�a��[��riD~/��|gě�T�S;5
��9�Vh���XnN�저�e.R�� ��'�-�i�٩ �E��hm%crN � n	Q�$9Jv���\ ��'��tp*��Z�x��L5p�v����~/��IL���ܡ_6*ژ$�ѻ���n�u_��Q�3���!�ߦ9"�y͚�1���UY��q5�op8�q�5)xL�y�Q�"/�q�#�qk��d�B�Y$L;A=(~T�X�-�l.^
v�2Qs�s���aR�l�@�3�$׹���#b��y'��Gj3瞥*���ߧ#b��D\ �65�^1LV�@ե��T��;��!a�~����aN�y��`N�i{�Q��_hAT�O�K�d31�fE��D'�蟫��#G�w9\q/ia�-|"2Ff��B��A��%Fs��v��h,C5���	��uK�m�p�&�s�ɵĔZ����i�W,�០K%��������HV&�Fś��#�����D�@��d�R�( �~}E�z$�s.��T�~T�2�� ����pjh����8$D�0��^^g �v�~�y����J6:��{Pd�.wK�6*Xs��tౌ�p������w��c�K����KsPע�B�������&X%n�r-�$x%Xn��b�i��]�����5���a��얪� Ȉ@�A���fh����u/��������փ����CϜ:V^�{��o�5�g����JF���=R���v+�I���D'm�"B��	=��\tw�k`�Fb�K�-�2�c+�牊:������3Ǟ�?�i�:�|���Ч�EIx06o/)�`σԘP�iaU++�3��5ݜ5���-��2�g�1v�ր��У�݉�j�*'J|9vv�
e�9�5�-/��́\���s�=��DA�m�	�����wOC���;����e�1�;�A�ދް]`I^��#g�n@����p�C.ŭ�#wAO1�s��]�5Ys�j�|���*��t����PL�nw�[��m�m�ly�T��;C���ό2|�{�Q�L��D��S~7�$�(�� �UƲ!��߇O��"�$����,(g�~��V�4͞�<� O�.�/Fh=��n�k��ϝnN��6��ϙH�[�m���9l+�'��,����H 4j�ȃ4����,o�8|ϼ����d�`1�6�D���[k�i����=�6H��s�1����'0�l��IT��V�Vr$�app�f��FzS��0
g�AF�����x����[�b
q��OH]��ک�5L8c�(�MǠ翩�����xIց���<m↎A"#�z�QO;�����G����H�B���֕�L^͆������:�<��p��rّK2�KA�&û�Ԅ
޵TN^�UR�i��\��RV��<�c���R��J���,H5��T��Zտt�&X��T8HԔ�U�RqLﱖ(��[�����e�z������Yrj^]��A�<Ψr L��w��xeo�T�<Bwվr��G�܇f46��GOa'hQ�����_�~������S���H�;.1[�(���ם9����wP�J�a�`��p����gs2�W����Ӷ���
L(�����l�4J��z����02$v�
���=@rv|>:ۇ�O��K�I_�,˧y49!��Cx�2�&7i�!zk	U����:��/��x�����qG��?��e��(�lدo87��9��˜'W�%��`C����B~	�X"�e���΋ ;�4Hd#Mr���r��H�OI;��L�S������m'�����˕���f���AmΜ�k��@i|��x��ۛD�:��T��.I��� �,�p]�ƪ2	�����b��Vz�9
�5���5h9*Q�1AoB���k0OДK�W�G|I��y:, 	Udpl��Q}�c�n��AB�(���j�z!�j�fў��sgq���@���R�:#ˍH��~!)I��*	%���|'��u����[���&�8K�A�$)F��q�Fq�2��	W�iG����ݛ,�O��P�������8=����[tK�Ԅ}e��Ʒjy_�#󎖪iUr,� �J����RÆ�3�R�t���ˁ�� ��v�c����!�a��n�O-/��`�g3�Z� 3c�g
�y��KV�ʖH8����!�A�)	�#�����B�/s��.��2'�M!�Jn��� �J�G+IZ!�r�b���/4*K����@�����|󼉏K�z��H��U�r��֒G��ٹ<�Y���@ 6W�W4�pZ�D��"�8-ay?�F�m�<'.b�RH��U��H�,kk���X�d5�4u�/�ӵp؞ٓg ���m��H�΋}
�����V��WrC��I����Xn#� ��w���3�^�#�Կ&������0����S�#��oE�.iq:��q�Hoo�Wܢr�D�T��jB�ځ��\X�Ś�Z��lP����Q6��-��?A���U��٧�k��^O�%��y�w�/���b��RZ2��4��j��2߃��3Pf�4��b
���ˈ��0��=�Fe���v{b��Ֆ&k&M<[<���ݲ��I�p�os��GL��%��:P���4$�� Y��Bѱl0`齚0�����9n �����*g�wn�2�\�룎�2�����y��x����V�8v�3����9�diW ��CJ�j<�N�p�����q(�y�n��~0��l�8�@�2����g�L��k: �O�";�U$��3��!��͚�����4��'�A�'S�T4�'
K����}B��ҝ~�f��o�,N C��ݸ&�]a����G���ֿ�<֙��8;ߍ)c����Np��:y��a�x�I3 ���-��lf��6�,��b�]+_���5Q�/�Y�w�F6���2h/#M��w��V���z�Ш�L�ݗ4ܦߝ�k��.ZK��K�~�j�:e� O]�[<LkW�]�L���l���Hʳ&��I�z�t�:s�^�=����>�B[߁��$�1�>���k�0`B�5���;�Il���wc,m\]���QNh��f�tӳ��?�;j/f�ܸa���fg��֓e.����:SLpeł祦���6�.LO�.�3�\�U �Znak:tcc��t��+���]B62�:��vg� ��8�´0�S�%��V �<[�S�ŕP�A(_���eJ��:]�Oq�ʺ:̫��Qx[1#��c�M6�����]��ӛ#�ĜbK-L�ѱP��/�w�Ϥ��~\��^�j����&�EX�e5����V��!�g���
������<��`����`��K@�$"Y�����6���^�N��$����`�[ |��T�X�����Y�|��dПɎO��{A�_ҹ��F���i�s%��J�ʣ�{���(kC����q̔}l�R���I�$1�O�-��
�)��%a�=I$w%��G@*�ހ�@h�#��\�@|�˺��(�u 1�|�hն ,���$���&�`�?�IM�M�^e���g�¶�j�RA�\���\���O?�7��P_16�+��s�n�6��\��g\��W�-��6��#�Ј���(��������ZpR^�*p�=t�/�Mheq�8J��p��^:	'�������pc5Nu��]�Zq@��Cn��ᒳ�`�\^C�k7fQb�a#���&6�Zi~�
3��\ǵ��5�(3�G5_'u�Y��G�l��q���^rŔ�/����~�<'�?@��CEL��/����5�5�$!����0�95�����?B�-j;K������9�;�N��I�2�����A��iIB�J< ۛf�w0��<u���F룓�뜦��uO��j��l�xԫ�r��(�-vc0�39���E�m2:�����M
�A4�W{��8��҄�:ջ(a�����?N�.�Ք>͘D۲*Zψ���;��~	�Ｌ~��X��kLt����(︔=�兤7�r'(�����o�M�rt�n��.���Aγ�"����|���i�T�����?J?%�E�84T��3�^m��j�>t�X��mh�ٝ:�31�Oܯf�u�ui}��hա��Id�[�:߹A��Џy�M߬�4�K9n	oITx]4�i^�f�5 [�[��pi�:�z�np�]��U��C�!Ȣ���y��l�P8N�y7H���:�Մy��+4f� �ƕ Rp��9��-V�(�P���B��!��졺�Aa����y4�$��r��9���Z_� �s���|a-b��:�<Fx{��È���>�qr�|����VPe��rxQl���'��,2^J�vV��]?���n#�g�U�c�1O�%��s��8un�ESgv�	I��s�Eh"�'��#�-�]"������Y`c@�	g� ���/]� ;T;�8��G�/�MM"�ڽ�����t��4/[�/Li5�}PiG��!���pg�A��v���v��),��Z�ˢYv����X�����4�iO?��M��e�O���ҍ��&����J��K�LL���3�V+r��M[w%�R�̣�	�4f^�ڞ�������gb�`��g���-�.Not���#�`���AtÞ�i/lߎ�{f�V���奮��	uݐP���P�C3�^Gwd��(�� F&���B���������%�h#��>|���Ƅ�����V�Ε����z�0;�P���ͷ����*2*}�G�{ P��<�g܅�vゴLN�ۏ" ��m
�E��C�_� ־��|�i��A �}e��m�Xm��p�s�˜�3L���נ�t۴;2,7��v��ɤ�w�h�,�<��V������� ���g :��z�{�>S�y�� ��R'Ą���#��3���J��L���4�(,�1oh^ѓ��3սŏٛ�����M��o
����SGnŲ�t���Tc�|]핆�bhfBI��]���ɴ�������B��S �W8�0tf��������C�����=�_?��H���F��J�Q}�����;a���ϔ������ɼN�vr�+�Z��	��vtik-�����n��8� Y*�b�lڳ���ٖ4�3�j/�����l�	�W�'�Q�7�c�N]ؿ�e?\y~��(��^3%Ќ���M��?W�����p�J��z�\��3�9��/mj+V�=�vb�8�o�d��v�v�Y���.���nP0+jʓA�<0<�.�T�h�����'�1���f�[����]R�4�/�D��_����/����9�^6��.��zCa;H޲�v����# �X�YP��{��0KxGy�W!�/�u��t�1|�B���口L���d���#���g�uD�Kӄ�+�͐Z���k��;�[Bξ׃;˟�.���j�}/Al��L�z�C،Ev��.rqʑijƄd*	 =H�53�O�V	���+���ܟ,��ı �x
\����|��1��y���Ǧ�6�s'�SU�.��R���$�E1��f1��޽�|sbLe]�؟0�3�+�IdMr�2v�y:��Rek1k�3�D{�TZ�/�LD��	h=�ק��E�b���K$-^�E�k������j�-�S�n�=[�ʲx�3t�.e�����Xv�Ϻ���AoZ��-�M--Q��w��Ȩ%��E��±��8A�b)�D���qo��|�:�@����:�O����,�Z1��>���p���/�Z����y5�	�ֈ�#����&\x橊�2ӮG��^�7OF�TI�3��թ�d����U�Rj`�uu=|����2i���Z_BnW�똡7���]�c~A�*>ņ�Nǥ>�2�p/՞K)��n49���4�[�Ե�Fj�3�\���FąP����Ļm�ϲ$w;��Y��ʣx+K���ښ~Cw��);D{��$�Ѿ�t���N�����
��h��BG��|�/N���A�ޮѨ-���2��0�r;��W1��x����7k`0���c�Y�`]��p���q2Vnxqc{�`^RO^,7�2�tD	As5?�I	b�ȧ�Y���]l�����2�k/���O�p���&o]��(��L�=hI< �iR�w�=�p�F����"��>�W�`{�؍?
[�#D�T?T!v|Ҝ9�'�T�%_�:z���*~3X~_���g�hZ�^���ie�@���7�$4�.���~�OGJ]xЎ��	 ��X��\��8/�*�2.�"�����^��c���Ш�L���I�8S�\��{2f_�{\;�.����Ie��C.�y��R5�nE(Wk��g��]���֜�}y[��P@�?r�xfz�7�����c��}wy��&Y���~9U#�+`����
�D�����,%�HL.���&f)x�.⬮�p��m��Ӥ6ydcJ�@iS��"��	-׊��-r)J`Ee����@0ha���;�mȵW$Q�ʫM9�4���E=�E�#$��Q�&+�c�e6���*f��T��]%uF��Sj��Ui`g����R���J�i~L߁K���Ocm�9������ԡ�#�䋒�\���!,�<�$���@����KMr�Q�f�s��V��zxť �#e]7��$O�0�ʯ�5��AJ������lP�
�4FƕQ�����M�Q?:��Ex���U�b�P��8�ܴA�8�r��I�H�x�hɋ�O�e��%��Q�<���TZ�l��Ğ�hYV5�B���dw�վGpu�����Z�A��h.��B��<��2��y��Y,f^�Z~���IA>g6m�l�����o��Ͼ�����~��>����Sun1��7@���:p�;<�k:���y?ifɱv&yI�VJ����d/$��;���^���n,;'W^��2����8�%���4�;Q���U_QEQy;�~W�0͹�č�c�{��ó��`��G�7Ќ5.�
bl����{����#�HB���NɄ��}�i����6��iE/��k�G�z�>�|Q�JqM*�=��(��!pp)��+V���T��Ud�1�ȿ�[_Л?*�цq}L��R���T�y]��l�r��g;��"����Q��Y겣>���T2;b(��P��l� �E�.���[������G��)pu+�+\�U9,L�9aӃ�(���ρ`���7ꀺK���+��4,���T�sF?L��Z�?Y�-���;[�#VxH������=X)�����o��]H;=�|�`�t�}���6��9�ɫ3���ʩ�#c-��+��,�0`]�<u�pB����v A�Kd�D���G�*D��� ڗ�+���_�Y��6����ρ^;`i.u-�����;��r��~k�7�w��=j�_P�*E�-e	��E��-�]��|��21M��4�"��NeP�N7���aR���iގ��YЁ�VRn~�"H'_z1�f4E�%]�X��2
��`�uX-A�����Τ���b����"��q���W��U�T��	�(���_��r]�n���l�sY��s��;�%޵Y��!�Z��;{����?{ ��&|~}�-hֵЭ����y�B�zW��;O��ު��9ț�}�6AZ��@�X��Kt�]��K+5Z����˭���_T�����a�P���ￖű��.�	�z$���2�
/#O���
���X��~
_���9�!:&�!��a��X��1��ޤt��tV,�b��_��Y#�O����wu������,���۪��\(�4�eg?����D�J������h�Li�QB�P�����ltM��W;�1�جL���\�oζV���2�Ɇw��qq� ��xΟՖ?Д6_�Y�� f�\w ^T{;)u�}1v-���K�����y-_Q�j���h�^����ȍ�8AX��a-���1Bd ��3�?�{6�Z�s���wU��3�#�����\��M�үI� 
�%9�H��#�Җ����ݫ�YOG+��z%/K$��.,�O�۴�o�Ɣ+L0 �QR]S��e(T��qaFB�}ԣ|<�e�v�ļ��H��R��%�f����a��J#Mt�.��S�ȩ��m'=��{މg���4#���w�*L��yw$(]%ŀT��-��Ɗ��ߋ� ҙ�҅�i�C�n6 ^ߨD�l������,/����x�3擃�<�փ��Cښ
>����x}��+�i���C�T����nKو2����� yԆ�p�B��x�N�� >��#\i��:�(�@0xC$�fj�4�c�7&:n��#L�A�j)o�P]�"�
 �C���Ѥ�dR�7g6b4��7pd�W��8�������y�g������ƈd](��#[!�,𙯔����]��K�4��m�`��S��~���(�+�9��c�?@F��i4̺(C�=5x�M�����N��'(�y��x�,4)ǌU=KK�Gf�G'5d���{�pmqㄠ�ԥ�����B������G�l�����8c ���S]�\{�?���Z��i>�����A�fW�Ŀ� |ǟ��ާ�����&,ʮ�)]�h+�LVԴ�U�pM�3Z'�AI8��,�k.)@��='b�EP���\ʗ�- <���}��u�|uHՔ���c����CV�˪F�@�4��/�:��	&%KG��lJaI~C��e�Oq�N�
�}CE�8@���smܗ������"TτӅ���0p�����ЇNH"��
X,�S=1�^�uCr0�y��j8G��'S�����:��H����r;�LG�88���?~��k1�q���.$O�!O�
�@�8e��`K8L����)��'屠˾)��?M��������R;t�`"FN$�I�]-$����H���#���֭ӔXJ�傒q����_���z���<#�aP�,��+�M� %�ѕ��$�%�j$6b�V����]#Aq�*ɘVuy�ϰ�>ZN��V����'�a�ȓ?��z�t�T�-��?C��|Ps�B�*<ŗ�4+S�o���[�K��8(M(g����\82�&�Q;?G��*��E�
D��̴WJ���������kA;��5�I�z.�|������$�h�q����Tg���o̗s>5�~��gRU�{�O���8�G���ȇ�%�KzRiɿȣ��>����L�?��
Sq���#">��z��AV����m�LY$�Tg-	��1��ؚ�R�� em��b����r}��l)��Z�b��\dZ�$�u�}xs��ep��0!�@��=���0�xroX	Yp��x�X@����EH?It7��/��h�z��|jz�P8�>�K��~bkk�p��q��x�������))�b���S�{k�]⬩o�
���=j�^�z�$��d��9������>�� �4����W1�@5��dkg��q��r�w�Fƴ"�d������W+���5O��|�*�`Z��B0�ȦZa:��?k��'r5�қ�*X�hy41o�D�b��,��5gQCTa�X[*�^�79CG�D<��a2��{^qr�緼�	P�ݭF!�|'�6�����\:��[��흧a};�*n.��}V��L���!E��e	JC�� �o?Ft+X��r��9^#D9���c}��*�3�Ǥ��E3X��D����xRD�>�;�,�K��,�L�D�~�w�=m=�;I6b�=��L�s��2�i�7�E& O��eft�U���,ci&������ܨ���{���B������	�	i��w�7��C�".���j-�#�2K�h0e��9r�;����w}��o!�?ϯ,�-,Amk<4�����"�AWcby�V�/�����(?��1�\�lF�PEX����p]o�{Hw)����
��8�A4���N3��#�4�E0�t#uSYy?����Ň��#����K8��_��gu������@�%Pܐ@��x����}�:-K�������;�>�;r�����3g7���BZ�ɂ���֫�+���֭�	���Q����Z�L�1�VhX�-�#�Y�÷�
��*��cvBj��fɹ7�l=��Z����)|��=�`�z���(�[�����ƕ���5��v 1r`a���.MԎ�t����ޥ��9"{j�5��]Y���u�r�^l3��^�w��,�8k�ڱ9��	�x�J|�	��A���Y-o�
�x$F/��`�����>c�.�SS1������'���pZ�S(j��w\�8������'��ƛh]�K%ߗ�0��1�ݾ���j}��D�1��<���CXO#��C��S��?�|T4w�B�0��� QXD�sl<I����Ÿ�,-�!W.EY��8E)ڼ6Y���+SG�۶ְ��`�|̧>��'d�����3�aw��Ek���ڴ��i^�|v1��L���Sj���8��QLSJz�[/�%0^���qLKe%�v�����ni�ű*��4�����i}y�h�`����k���Z+pM
iJ�F�"qû��V��+��������,�gB��l/ �9#jB�[C�,p6�*�^��gQ�N�9#V�!*()+-�����ڎ2 Ap�N���_�������Tg�N����8��6q\*�I�Y�;�������� &&=n5Ƨ7�"T��Hј�緷]0�+Ϋx����B�q	�w+����&��W.y�i�:��t*�K���q%�j�����VU�Q4i�%l��u�3J��6���h����;�96�J��I`��aG�"��|!_8/,0����m;���wu�Х��;����y;̵�E� �\ꂍ�)�u�M 18I�`�s��ʑ6G��J�N�8X��!^�dO�ax�a��t�	0٪����Q$��P�ش��G�iu���5|��9hZM#�[��( ��bADW���,ԛ�����[B��b:�/�H���Bނ��ٺf҃�ɢ��*Ru�g����� ��Z.�g�"��@x>�
M�B�[�ya[�*:s��	P�>��/�,���/���j�/_��=ĳ.GmNB�h�ٞ&�B��C��8V-O���s�&x��~����~x���n��n�ŋ�6n�|؂�R�d�K <��C�V*!�����E���?���ߴ�[��<���5�z���L�Q�֜1`Aq�X����K���H���C�2��G�C���ьʹ�`����c2��1���.����a4��4VEwz�eTe�!����|%�s��	��:_baҽ����J䳾h��+��N�������Q��Bl�Ҍc�hR�.�����O|���4/	i5S
j����J�}W�1y���zA����^�@���%2�҈�/���y[��~����VYic@6T��؆�P���
�
K����KQ8��PrI������	��&��_��~�UAF��Ak�/�#qI��N�x�<�1�@�f�*��l��Y)��?lJ��쇂�V�e��^�E���m(�,Ikb0��'d����d1����si�ס�Utz���1u��=5@*�y��i�b���$@��VR1�aY����9�� YQ�9�t�Ɗ���'�U��RAzJۓv��:*����ՑfN}�4�!��1��m'}e@YR\�L��M��=a���V�G(��5���
�J��-:{#B����ek�YP��r��?^EU� �'�?�kI�|Z@�f�2�D�8a,����M����
��FR�?�y����RC��A3�x��},��&]�{��.�7�_�2����=��IAU$ԛi�-ҀW��Kղ� ?��e�'|u��C����dY&	��>#��.�A�������;Q-CiP�j<���������CT��A����v03R��mh�j)�t���+uu
��%���N�����Z�<H���;n����m#+EGd�g�`�\�qq��>�s�K�`N5�l����G�,~�բ��v�)�֒ǌ�rpB�a�ӂ�yW���ڽyF�����c[x��I#�(��<1z�-]�;n��j�ws�wZ[��"���?�t"�+]��1J=_g����
�ı�wt�liʶ i�IM���ʃ��E-L${����v�{	�zb�l6?�č�&V=��O�e�j�َ֘2�0�T�F\����~x.���!3]Hϛ��I*��S��R��G�پ1���r]�����m =U��4kx�W ���K�<\���|����S��Vz{Y,5�23Z��2V ����K�{���+e!>��p2�x�hOe�clF]�e�Z/&�	��|�y�`����e��z�:�=n`h����&�
�ud�`�j��۪.�,"R#�z� �:�j�9��<�A=@|�Ǩ[}5�4d��IׁϢ+;�i�j:٬<�{������*�D�4���gr�C�H5�CYVw3É:��
����˔�_�.L����&~<a��q�~Q���nؐvb��ŉ��f�{��>� ��*cz6`y�6U���^��n}���C�/��(u���{K���U �����G�/[�0D���᥹�p�GL5$ ��g.���K��|�9��
�P�ݐo������u���+2�c�f?�M�ˉ�+�oE���a%�D�N�6�ؘ�mt{(��C���3�J,��/~i?ǎ���`}3J[*�U�f������?_�n���a�P�;��xv�Zۥm`����x��/�T�c�V�TpW��F��R��<�Yy�炝$;��.5~.���e�>���c:�.�I
Z@C���	p�A�0��7�n�Hq�>Qk�EqH�nM��s�G|��(�������/�3W|~m�}Ԓ�Q��MAa���P�h��aL)��� j���y����gB�F��bX�J�O��t�Z��gI��]����YN���B��	gO@mp`� c�z�����I#�z������K�I��YbBp�f�bfI��ӟ+黕��C����1w� ����Z�R���w��'��D�V [�-]2��a)N׀����b��Ky�Ͳa��'@Ns�iYr���ʣt`"�����vlN��;�e����NY<�(�-y(qS�ʬ#��$��W�x�]ڀٝ
�z7�΋P��	�~���ܝ���~��
U����1�[z�����9�*������Jr�f�>H��eR����(����bCa�}���R�@!-� �a��la�ٽ���:���a��G.I��$�S]�1�_xeu���|����G,�I�=<�`i|�xy �XI��Op ��!���'{(ȊL��"�S����j�*-�U��&>��iJ'b��;]�����;��;�QOry��}��Z"��������D$h<��V4ؒR'!���������S@�*I���=�j��:�FH���=~w"=�#��"lj���.�k_���e�v���%0�J�;�K�?�cY��@LY����ezk��(r��TIfi� ��na�̹�͙�F�`�+���\�¡��r����r�G���RUh�
�)�2�5l��}�%0	
V�XP(~C�y�fT�O7Z_ɔ����� A�zrt�d{r���Ap-<���HnMP��,4x�|���MA��@�ֱ��,m��JR����|]�2�j�rP̌�|2FB1�pw�ڟ�T�dZ~-4a��0dڐJ��;_�����>�#�^��Y��NI��a�fƮ^��T1#R���
�k1�ĥ���Y����#���Ĵ'�Rѿ��L=a-�ө���q���5R
Gfw�ÜZ���z��8�l�� V{�,@�zhӜ��X�.&���+��pa����9`��}�P�i��lk���R����W h�~�)�R�AFl����ב��X�4�v��.����D������@^7v���qPs���E��A��3���#�aq�A��?��	�h@	3�>����p�����fF�uGV�,ւ��pw^���E)1=tU��Ĭ��:u�a�d'�B}o�?�܃��_�u���K~��/&m��M�I�-|<�ԤO���c��B��Wbm��FN4!�
�>�;H�M�j�P��U�p!#3���x�`���Q���L�,S ��f�5���2�0�����QM�M�Sr=j�퐛aF����pYCx��	E���o0�p��JL�i�9�]��ˋ�4d�_�}�&��i��イ���l�Mp�q�oc�,"'��I~��A�Y ���Y�64�����Pp����:)�A�<�osp��U�-��z�xB@��%�񃣹�+�B�V5ւ?�!���Ht\M��:����2_�s�9�A����N�3�>���{��3�p����%/?�J��n̳���e-�܁�83�2��%���L i����,R�i�$��l�z���,wR[�jīV����qp�����1U��Zˣ�@��P��vj��������~*be/��QK��-ɜ'rϘd�v蟵��4��1Pt�����o��e��R��/7�L����P����q;y��k�Q�KΏ���~��i^�D�li~Y�\D���^�P��)C0�@/g�	9�@`��z�m��D��sLJ6��X���#U���q̛�R/J|
��xh!
��������/c�=*q���+�4/�:��7���h����� �Mylu��O9��C�Q�q�����f�v|��P�+Kp���C?��Y�\71�~U
�/=��5��Y� J�wVx�RI讝���Q:��>�G 㜬 ����L�}qǵ��'rH��өtE�wC٩��ζ	��.���pG��;��*���%�b"�-��`�O+�e�J�?q��j"6Z�k��=������D�V���0Q��h�a��j0xl��]J�	�1�j�|j������GQX�e+�����~%k�E��}L��#�UD^Y�3�7�=�w��.Yyn�4(�T錾~�S��Z�i�U0����������Y i��Gs���=F����Q\�u���1IϞ�I�o�2�/��n=~�$��Ĭ��o� ��%ŗͭ<�o��pY�V/�m�kϐ̈#d0}I^�A"x�D˿��ǳ����:�Eqd�C��%��.��I����c��ED�Uhr5�ܴ��Ą��Gl�b����o��[=����8��#��w�h5ST�3�%�O��*U�h�uz+�+X��fGD����G3m���4}r��ܦ:��H�v��@^�P b9��
�g����(Y���%��u����3��HlVt��]�!7R��C6#$�EJH��:��N�}{[�%��)r�^WEx#�e@:��Dy���!.yt�p��'6��%�.	^�FN�+'-�혮��v�L�	9�W�% �K�-k���PΎ���:<-� B�K����-ֳ��"��t<S������J�h�ł�4 .;���b�P'���z_�����P�5q��5{�0�C���P,�	�M��R�T �_��y���`�wTj�.3��o�d��ϔ;e���cCmyЃ 5Ӿf�-��������
�­I|��U��y���x3�u�e�̿!3��5�!�#���Jd���m�a;y�/h�~��PW��1���N��U�띭fx��nN`N�b'Y��H}��	�X���.��*m���\��鰩���d�	K��#6~*��@�T,�x2�
g�D�SmF�}�ov�)�T�/�7�G��E�~]�3�j?9�d��A�|ГF����C���|Hu9L��]�!0�v�2��D��F�$�N!7f�h��4xۢX>�y���8��&�����§��Ĳ#�V��Y��11�?A{J�Y�����Ȯ2q]�a.�6j ��\���)�Q)��_��mA�P�Z<��� +���ddL�sԚ�ޮP�о��n���������!���]T��m�:RV��;o��`fk��k�ث���kt��wp�+*�5a�Y�d�F���b��p��&o����ЩLC3�f(�r���n�� ���R@�?�(
:E�����|恃�9$6�8�,F�e��:.(��_��m��P���EH$�w��Y�1$p_�+GҔ�وD*�:7�h�i���N�3�[�z+��o�ξ]������B�Ԍ��p��('�>���Jv
�Ʊ1A1p,m¸�}��6��諒`�C%O6xO����O�����c
�� Y�2u�����|ؾp>� 0c�q�\B�Pk�#�����Y���rP)��{�o�v{�ah����{��Դ��cgS�MmM�� �Y�-e� m8�9n��WXc������7Dx�q(��0��ϤߡOX@�IuG�86�Y;@���1�M7n��twxʃcB���
V:s�;���M�R�����[����C69�7'�!'������ �}���q�}/��+I~U0�di5W�3�f8�1�"���&�ו�ϖ0kj���])�ڸY	�VF)��۾�n=m9�M+;�g�4�h�����m�_�^��+ܱ�ڂ���A��"�Tki}х	eɶ�+�h8�I4b�-����8�]i���)���11���͢2A��3v�#�l_�@p�m��p�D֠v�3k���>��;���(��^������E��������O��C����;���h�Aօ.�[�"���ř	�p���Zd��~؃)L谚{ZҪ�H�*�&��+�?^:����<��Ii�c5�q��U���c���X���)�H�sK�!6��s0�i_�jV��4S��g���8��]��U��M�������+�#��n�S��+�jxg�ְ�k�7��(b+�h֜x�\��3,'I��?C��Z^Fwv�ao�{�((��fe�{�*���E(���L�W�V�c����{q;ݵ��n�.+��`��<%>���>�j/�y����&� ���.���=��/�i����2��B�L�߰�U�����+Sބ��:�*Aq˳4=1T&d=ց�T=ƤCg��u w�~ގKI�輩FK>S6,��Ɲ�Ui�f��}��z�}qviኽ<2�)�aΰ�ɿ�Z�L���2����� �r-������6�W��I?z�)x��X���DM����5������f�t���;�"��a�k�ga�"�L�ع��~IC�+����kG�8K��QxWe�H��������AZ���Y�jM���"����[�sX��� 5 {x9�V���-y��\�:�}�~�g>e������ͧ���w��)���yq
	^xE�23ia�5F�3؞ԍ!���tȤ�y�����5Z�b'�őT��a/�݋9�����w��	�(�2����m��B��x���'��gƒ�s{��5@��D6�:T�B�N=.g<hc����+���۰&D��@��l-J��ԡJ]��}�.�*�j����������B�]iQ��v)5�UR����e�T^{�T�B�Y����&�}@����X%V��݂
�����e��̏�"M���21�Q��6O�K�H�&h�d��qM�CU&z���h�6ߦ��WTLLMb%�m����J&��|Y��1���fC�"�����Y$�� R
PLW?Wڳ���\&}z�4�6�滆��ճ��d_�hׇ[~��w���(m-��{4��o���[�nKv|Io 9#^��=IFfr�x���)��G7L*����R�Kx`�����o�łܝ�(HtL���#�֊��y�= �)�L��'��Dν����(-��SU�q]mIe��8t�\B RM��;'�s�m�ɂ��K]�ۥ��u�� �zha��Euc���#��3De�yt�*6}+ޏ!�Y�C�cM�]���$��S$ZxZ�B�ur먞e�`���<��3�f8�<��_8C��T��0�W�n��?{Nh,浻��d�S��_}�ʍ7��T�\T�����C�����ݶ;�Ҩq�+�^糰T��mxu��.��#���FE��+L&�m�z��PI����ϨH<v w�o>�W���d�Uo'�@��}���QH$����1��� vM*]��gf�?m�A��5�t�`FzFV�A�yu;7�L�e5
����G#� �*��~X ��(���N�!��rS��I�����_
:����ˢҏ&U���/*x��e�Dр:GBT>`�����Vq�h�1�|��z�47M�m�m��r�+�/�1ޞ�c5�T�ˇ~�+%�~τ?�L���](\B��������N���3����9��w��6�Vg�6�v�Cx3����dp��I���+1GS�JӪ�_$�g���s��:�Q��i�^R�oM��/�!�᪉݀Y�ykɀ�R�ߦ�/#`�����*i"58p$�h�k(�J�:�ܷ���bx�B��i�52��h1�R�Ч'��tYh�>�˧6
ɣ'bi����\c75L���J}1䠃N>��&�ږǡ��;�s2�=H1��vԍ�Y@(��׀7m�n�S�C� ��ܤ9r���;:�-=C�?�!�>�0����<ل�0]�x��?����*�Ǳk����QfwA������..Oʟ:͑/��'n�	=��rW
(=�nZ���2���6"��3�ag�?�H�W�_*F�?*�������ؓ�m��:v"�}?
���%�>?5�*U{D��k-H���mY��mf�k)P�h�_?�_w�C�Ȓ����nk�4��L`\����]�?��E� )� $�K0����4��8����7���&a�n���ό�.!>=�&�>6ɶ�Ҽ�zX��c����&��;��}6��j�O��0���mE~$�?jm��(��Ƿ�Z���8�)�k�i�5���r�;�xDͽ�ا������_��ɧ����c�Q�)J�G�e����鏀Խ7�Y��r��������6f�/�j��(�P��t���?dVu]�8��k0�,˦�c+B.'3��m�)]#U ƛ��=><�xS�?�:-%8	��CX9���uC��&ZA���6�RQp=l�ص56�}	�ڈM>��k�|%b��&
���1T;5�dD��B�oTP���8���e���H�B�&�x��`����j<�7F���A>�;�#l�����\ze�*@�0n�6����fF��Z�d�A�j
�"	��8	�&�8��A��uc���wh֍�M��t8M�6�&88?�A�@<�XȎYɩ���5�rlhkL����#C��� ����.8%�Yĥ���`��j�(��%�G6���D�1��v�c�g���Z���Z��	j�~t�,�w^�gx�٪q|Nm�ѽQU��i��N��t�.ht�&��U����J�	:��Y��x�'�Qe9q����NC���e՘W�kA��g	mzlY����pb� Hӈh���w�j�>i�(������V�b*+�rF��E�V���i�g�.JY>�9��M�K ���r���v�"� 	;?r￀u��Z�ǚ�V ���ڝ;*O~�C���R#%$ k��g��z[��n�I'�����ʼl��l>�
|����;���Æ�
U7�-���EP�6K#�޲�g߷��o7ݩ���_�a��D�k�+n���$c�+0�-���1�=����QO�kJS�W�u�"E�C���l(�[`�3h����%uT?���fP������ȫ�����'��ރ#4��"����k���-z��`]�s�#��R�-�������$�"��0����i�Vy�����q���j}
��ȑ4i�ʏ�:�Ǜ$�0��j/����新�:�i�)�\	bZ���͜,�O�
7홃8��tH�P}�ɮ1�.�u&�V���C���b�);Ԍ���,�0*����L��z*�-C8�7w39�Ż�=�6����		Vfbmk�4�c+B��8�Fݟ*,�����j�'Y��a)y���(�����/����Ll6�H��{ ��O�5����\`w�g�y��S+}0��H��Sj�� 3k�-	�"�(�S�f��g�*)�)�>������%��}�f��}I�M����R��)��Ad����n��[Ո2Y��(=�NCz)˰�dQ��ᗏ�|22%��Mf�F�ɂ+���j�xIxv�y�e�495˕��f]��gp(�B�C� ����B�U\�IUtO�Q�#"��� a@f��l���A���^���w������I:fo�	�22y�pR<�cZ�q�Vv��,gD��g�5�֩��isȆ��{�󛝣������LI���:��@Zc��
���bY�@з?��g$�P�����Ӎ5�=sU@�/V6t#^��|�ƍ�;��#�9���Zԩ��Q�I���v�|Z���������9G�`��V����3Z�q��?�l@���뀈u�dm�4/�d�)��� 'v�~C_��Y�al��~|�RxF�f�]Ȥu����ı`zwдZ�aN��j�'�A�o�L9����:$�(�k�u�:���&<<!�A�QkF��r$���Jbk�G�5��XT�^�<&�=��� `F�^_uߣ:~����7�����ȩ���4��&.I��d�\�Whm-F��-ML퍧Fj�B)�^�%:� ;c�.��7h�M����EzQ�3�S�ƕ�8�R�T����3V'�p>|�Ns�; }��=�6{fe��2����FO�|�Q�Q.��Cŝ7� ��|��=7�g�&��Z�ҝ�Q��A�[O?⊫�/�s�`e.�������?��I7툾�:ٱb��3�
�ΧIU��R��,�B!�ۥQII�8��O�L&�c;�pI�=F�MQ�1��D3�ۻ�d�#��0��A9���\�7oq��
[9$��#���dգ�����&�F6IW���>{Q&�Ⱗ,Uz�7��l�w(�^]}���t���}�P$JfEe��ˇ9�KV�~�|Oy:�lZP�ᶣX����vY��ms�k�{����������DD���r�S����2�>_��9L����f�*�Dnݍo\��V�Ws�Տ<�\7���J�_��Ǜ3
�쾝"�Π��<��g�c��Hx�6�bϲ�rd�b"�O i�x�1i�8���> S,��@˯>�\SX,'X�J5�Mli�H;K�l��ι�VC|�`�Gt�#v%���9�>�VG�֖�zߌ�5p$'d�@�}�-qp��w�ٟ�:1%��p��#�)�>�:�I1��������5T�����!׏�4�V'�NL���1�n0`�.����ـ��<x�����J����OW�bh�J��[-�L���t�����ث,�/��ΜX���j.�y�iK�0R�"�M����_�Z�(`�jv���x�2Fv�	^.�B�#��(�.(mQ�>��禈W(�,����~+��}iOL�B*(�Cf�����|���턘��կ��������+3j7��{�I�a�b��:mzI�_��~�(�g��=���P¬�ȴ7�>�>H��j~���\ ���e4"dŀ��焨�kЉǪ݆zoÑm�۸��tF"�{�8?���
��Zj����Ԅ\g�DkF�ǫc���?���K���Pܰ*�m@�CR8�jq��첿qA��j_�aO��@�J�n�&�+ww�W���(�s�0�J������o@-W@Xn�~b�ptH	���T>F	:��e_����Nc��0���-߈
��˰�뒓��%K����^�V�7����B,��QWMֱ��;om� �ޣ�v��t�fB���=�i0����.��-;z�yL�4~J�a�:�-�T�u����k�N�MYn��ȤXwx'z�A����	���D��?�@Ջ���'����Ⴢ5J�U.��|��۴�5�����`X��T�@l��+lܽD&�$M�E����ǶjՂA^��:�EP�h�������������u�j����U�&�^j* P�CW]��(�a���w�E�J�J9����J��G�S�z��QLKY��m�F�n��{ƯA}V�?�_�6&��ד��Z��PIU�ư{��#��=�T|���g�$A0/��J�s�曯�BK���Ȟ����U!��y�-��'���o��x� P]P#�=�˸���$-�7z�7���i�{M.=��z����&��AMd���H�Y���~[MNĿ��~U��5�����9������m70c ֈ�u�y���̜�n��ae�7�J]W�*�R�o���nD�
[�g��CZ~���-�PP�o���8"c�`,��$�au)�ڻ��b�υ�on��*��ނ����E7�� K��E�]4��Q�o����^����4h\r��9�ӹs�jq;�!u�b9�|d5Z���/�`�S�Y%����щ��5�����l���d��h���َ,�u���{��1#♳�ف]e10!�"�Ӻ����l��З��a�9��J-=D�Ww7��ͮ2D�1=�tl���+_��uc��pj�5�*�玭��@m��22�ܼ`�I?~uMTZa�Wϛo#��M�xj7L�قJ���Ù�O���3 $*!~�j㔅�}Z[3�u٬y�Hl�+�p��aހ��*<��\/{E� ���U䗝�gdX�xA�t�`S������/'޵^��4]D|����W�4��������1k���Hӵ$��c93�1�-k��ԟ�)q8^ ����_�w����XUFD���e�%
���*�5ɪsF�C��bHv���2�#����V}�8�/�� ��7b��>2�Pr���_Qv���D���@��P��!d;��w��wDc�2v�9���V�^`K�\�cjԌ�L��S�ԯy���^�ݰ�bzI5I���׈�YM%�_��>
�0��Mg�L�v�9[�jEl�M�CG����x,._zmx�.�F��QT���������@��[��<|m�F�b�#>6������6���|�t uV�(9�9�\'/�h
�R��ؼ׀�3$!���NW�?mT�{A�]�c��ᅧ)��_�f�ĔuzQ��M�ߍ-=�����S�=�GNF1�K��x�_MK�C�0ɶEߟ
,���ݔ3Tvǧy�fv�e�&UTcf�e�@ʔ�V\ٗJ�Q������^ԃ�:	S�����⬥L�-�p�����+E�Il&y ��tJ���/%㪇m��4�?>��F��=���s�ÅxS"7���ޞ��� M"�\[���zv��C�(E�����+/޶�&d�PjM�I&"L��[|G�C�ax@-�K�OoJ�D5u@ս��L�R��_���j���R�����m�-��n���Q��y����g�s�W���|�Ǎjo��0֚��:*�18I�����87����
�A�-�����.@�HV.��(��fFi�\�7��#S��tr�I����w;_��l�=��ڏGTgs�w�����fu���GE��9���~s֣2~�W��:�m��9� [T���r��g��tE��l�00��b�Y�d���n� �7W�+�*=άw?k >��)x&̚ڒ/����~Tڤ��*r�O0j�D;��όgG3�z�H���J����2�7�����AX��f�[g4�Y��eU��ۂ1C���,76���p�{����J�}���PE
Z��@H�Pr�4��:d�aWB���Sc�@D��U~"���m>��fV�F�������aF9��YO
j	��g�Мc4�?�Z0l �s�S�>g%����3zb�|�a��)�K�.$ɥ5]�^R��F8#��,	�M�/�+������8!��N�:
�%�g �}��A��֪{���T��j#����Վsۓ��u4�GAO~���
�w�5Vi�v��<R]�
?kS�V��ePA�X��	1M`�$"tldY�'���f�uߧ��Bx8��`�u\�n�͸-	��ϕ53���J�+���}A<�-.`�����x��Z�����]2v8E�JP/�XO��c��5��5��A����Xi��d��(ϰ���٧�$@x��h���c�u%�X�	"��k�.�I�R2I��_w�-���c��.2|���<�pAc��a��X"�@��B	�xqF� `�!�n�ؗ+�R+���� ������#�8Gt�lsr!s6ٹ��֧�	M��߲�?�."x������&��M�?\�Zca^D�����~�����~3����]��RU�O�����ʵ���*�c�U7c0l�.%&.�;O,@�o����J���>��k�����v޴@�W�Ь��y.wZh���U�
�ώ`�x�����wj!p�4�Z�
^\����m.Y�� :X���B��l��q*�X���U\7��uk^���߿��W`���#�I�lV��XN�����#���gQ��J�ll���U�eMHҏ���� J�]���'�ٮ�Q��5�u���>�nN��؄��^�8��.����$aiBG>'���]+!Y���������h�Y7�|�1n�k�P=��3#�ה?�ꛪk�RF{p�n' Ck�m���i��kw���2�����D�'�}�$�ŵ���T��O*���,�^���*h��EI�C0#�o�-��b��\�nި���|FS�k=������2�����C>`I�B��Fu9��T��I�:��-p��(B�3�E[J�g&�����4������!�p��u�?�C����L��<�^�{�^�-}8PK��$�/Q�@��XZ)1�HFV\7ZRpxڗ�!���34X��~����g�w����ɚ?t�:��1��ڝ ��� ��!�7Qǹ��^z��}�+�jd��*P��s�7^;Q��j�|R�C�'��I#PC$e�
�;�o���]İ�h�m����Sq��6�<ڢ��9��.F�aQ8�V)�N;�4/�p�Nb-��x��^�xK��>�n���H)�����yd�Y���T#H�DK�Xu�����zG`0Sn���}a���ƓW;��**�=eqy���_>W}���Z�"�V�o�,2ikPU��挒�C�wA��ڢnRx��B"a�}a V�s� �Ƅ@���N�C�YAC�e���h�o���;w���M&uX%�p��A�]���cW�4e�� �Ϲ����M�"	���C��$ӛh6�$�]˻����:7���7�Mō�j��O_�R{@	��b���){9��%Ah�GN�rz��$sw��o'�O�\��G6���Tq��PM�S"j��-c?�+d:/�;;��"M��Ȳ^�.p_�'(og���?w7#q{L��g0�5�e�5"�nKgÅy�T�	��>iA��m"�2oނ�u]йp?.6�;����Ŝ�46NTV(2�)�3E� q<�*]C3�� |�����U�]����a������O_����c��VR��lM�
7$�[ƍ<9s�,�7��R��?"Ol��ǟ�]vz��T�5��E�j+����D�h8bS+F��$u6��'�	t��f��S#���:��5�Q�_Ih�#�t�>�6$r��d12���})?[���r*�nc��D�nT�m�C��V�1^�F���Ib@-��~^����r�{e�60���⿟��ue�jo���6��#�n�M��~RX��zm��~b�y�2���X=�.0����~�z/�;�۵�CzX%��6���2|�)M�A��}ژ��������؉Sn���C�%:�Ljc�}�qk~���ca���P�^W���w���z�UP��&C�*�2(� e�LX�`o\E��I�����8�8E~Z)�%ii��BL��*16)�&P#q���������<g-�$u�-6���U�2=����"��.���D=⮧����Ư��2�һ=�$��R�;w�]g����g]�q|uG ��L�L�!��ژ��[Vx/Kq��?�\�}�(ۑ9��7�W�O�R~k�>C�� _�l�6����٭֠프�䣖4ӏ�����i�Ӆ�`�X<?@�/�@�{3㰬��5����X^іw�O])Std8s@�u
���f����!R"���8N�F�$?��h{��	��ꁲP�q�Y�]�C.�q�	�y��*��4+B����+���, �]�N��Ih.����#V�F�{Z$�93)]V~�_�XR�,��o2�.��o�5ˑ\��c��!s+�gofp*��sW���\,X'%����ot��=�sKN(���R����$�G6���[�J)�i��uܣ���se�o���Gk�� �gu�~n�ß^�:��c���&b <�R�*��Rb��;� P���Ki	}a>~����^�a�X�Ǯ�
�ǿj����̷u��;��N��R�+ik�"�~~*��<Ojh��:w<ԎQ����0��.��,t=MX��$ W<lt�\�5��$R���8��]�����@�Sq� ����t�o�Q#iְ�Z��D�g��b{'!�=�l(K6����c��g��i-��S7q>�o��ʹg҆��~��F��'�'^�M����bS��!@����x��p+\>�^�!?A�Z���aX���m�͖^>q��h��q��xhK���M���ڨFs�3(j'�4l�Z95�D;�!�xD�,��~���4;�������9���|���&�كQ�Z�Dz���^��5�� ��AJ�W@�~�XP����Wuc�f�1��KT���T�h��L������S�Bf�/+i��[�q�\��1����$l��n��|.�P���mSϲ? |�߯a٧��yq��&D�����F�*n�"֟QTP�� ��f鴱R�u|Ŋ.M�s�Ɋ�(�����l�a�מ<��|$�4���,�K�{^	�	�v�$���%/�CC�}�3�#�}Z���񈺜��'��n��C�tԟ�9�����l:J鬌CGȧ��BIo[�p r�OR��>{ʅ�#[C��$�C4X�3��D��O��i䜩�qE�����IY�Q�N.EF��$�s�J��`٢���m��RVV��Υ�D:�9�
�q��*�!!>���3W�H�O��֭����s*��e��+`�cս���q�Ix�B���]y��靪��yPw� ��ծ&��sQ���k�c:�_2�n�
�?,�mtp��e��� 1�y��/���@:PJ�`�n ^�L��u�5�3
�G ��3A��h(���л��?��g咹b����2n�Mx�p��]��څb�O\�gB�f�r%g�'��DU����K��7��Dύ�Q];��?����e�Xؒ�������*�t�͍Sh�3�a˓���Q�Ead�M;�<A�R�hȬ��]�Z*^3=�0�ʂa�刻���S^��l��)�stK���B�"`�<�]����J�";����4�J�.��6"�1�k����y�<~A4�� ^�2�
t�4���3��j��2�.0��\���
�2��ҳ�5�}*iZ����m�o�9�v ^��G�JJ��㈇�e4h�.��ڋ����.M����8�Z����uI*� t%���^t������-}D5`q<~]��(ָ�^2�c��E��%�S6Jo%���oj�'�r]>�S&d8�ϵ�	eO�ʗf������ם�O۪��i�8�
��ބ_�C[f�q��U课,~���T�sWQY|.DiD7�_�@f��f��ր�Q�@.޳��I�N9��9c'�����G�QI�m�������ڞl����:�(;�1�Y�M�#:�m]������%���WpeS5ʣ�;9M��7��R��� J���M?Tfܨ���l¾@�Wt\�q}lLM�6xv�7Ŧ*���D�&���aRR#dE�Y��O:�ֹ4t��e��>�.r���KF3�,��T���M\�% �)�{�j����wAv�,���:�:�l,��fJ�#ō��n��ßI`	�3+\fխ�������`�+���Tc�;Q9͗hn~�Yt(6�Z!Ec����Ⴗ����,#���|w|[l�����T9W������j�4���z"��B��9�y�hR�y�����f��-(��v�kKhr�)s1��y�5wݧu�K* n��Я�+ZV�ed-&�툧p6�''�SyI� e�O�t��M��%�	�)�h&}a�-f�Ew����c����8Bh�[n�B�Nm�A�H������G��Ӟ�/\v�t������� �eR���s,thx��{f�4#Q^�S��~m���Ѭ�{�&�GF6��xRQ`�A�7a��g������*��x`��~��g�ʷ��k������#6|�N�n;R+�����/K�s(P�Ѫ����R
U�U�q���
�֛�d�VJ�-7���0����O��'�Z�E[8U���,KDM1��yiͫS=��T13'	�X��y�fB�S�d�8b��_�������T��Yaݡ��}�M��N���^(u{`D�Aw�<�v�r��$���Ȓ��/a�AiB쌗M��O�0`C��Le
9����ωD�����R���0���N���g��ߚ�3�Jgӛ�'��0F��7 �?�g� 8y��9����$S+��A+Y2\K�u��<)פ�w�w~A͟�Q��g�
�c:�0��L��7��U����(b� ���V��������ŶP���*��Cx���ʛb�����A���/1��jr���ɳ!�&Pf!Z0oA�_9���(��BՏ<���-�P��,Ǖ�K�8_1d���J�Яg⩖�_-������s�I�5�X/�*x���gt��'%�z�6�R2���o'��#�X�X !�����$� �S�.�!y���
����*�6I�sC`��wlC�&ޢ����T)���Hۺi�oǂ�6~|�5_Ai
�Tv�4@���Q<��x��3|O
���5.>��+�k���5���lg�M�zG�z��d�Ж�y��������Y3��+KnZgt���[$���x�!D��s�j�gȁ�_b��.��W/eI�����_Ĥ0TmҞ馊�σi��Th|`�Q�|��8_�RC\<y�F��I����5~������170��p��)��:��wdݷ�B*��u�L��#.�)^�^�����������؛�?܁�����_G��m�R�35>T.lv�(M� 4ؗU�{��F�*!I��,}�)�}�[Q���"��R;kl'��T���������vH@�a�8��W��b�\�r��f	ӰN9�^(���㖌J�Jo�s[�\�e^���ǖ�%Mk�,TL��B`u����T��0���B��mzu�
�(��O�0yQ|���i=�0h|8��M&c�QXV��^7Hbف�Ņ[}��i46�uB���W���G�$Z�ρ�r䜀Q�|ޑ�<�C:�6�F��O9y,���QH��S� Zw��m7g���R���]��5#��BINW��+4���'�ލ9�[�&�p[&��{�&-���h��!jˏJ��x�Gu�nb�d+�u^�8:L�Q^9�A�&H�0���rE��lg_�hj�����ߑ�	n���Y�uv[h��반�%2m���FsRjrW���������o�B!c����=^���5j�dp�0���
]���r�ɚ�V�������	�Vb��D��`�E%�3& ϥmG9M�uգ�=�?n���z����������@NFF�������P�K�Rl�1C_G�v�G���BJ��b�6)��%߲#A��9����H��4Z�Y��K���|����^�v�q`�`9IjE���z@`h�����ۮ�c�AH�c�*R��a\q�+��A�U-�1�&Ғg���C���XI����-�����{� �:���GԽ��&�.]����d �.Y��X1V�v�Oӊ9D9��&���(�T����1VAxTL�@�l�J��)�rM�R����	�Qss��(�Ƅ#� UY}B�NuB#��:���:�}5��fl�B���ϔ�����N�ŴC9q�~�]���-����� �����n2��ʁ�[02j��1��J���f.帻� 8]{�Oa���6�W�_U<����ԥP��M�*�<�e���������(\���)�1�B_6Y�b��T�o]S�!։��>�����
���X7i����ѿ�����zJo�_Te<PGИ^�g$ӄ+�q����6P@�|�ë�
��Y�7ً����i������n�����N��x�+�s����]��`J�+O���G�\IM��Ik*�~��wl���R��E��:p����r*ӋQ��/�q(B�x�R?��{1��X��3��{��X���Ŋ綸�]bS�6Oͅۃ�~����LHt��[=�{��M �{j���u]��&#݉�Eޯ�Nw�/�*����z���y����g<�)��LM_�wp�u|�7�b_|�z��XQ.T&Y�Y���Y�D�QC,.���Y$�.���50������ֆ$�5c�%R1BP�Q�)�*�^bS47�D�f�ø�����G��+5���_H��-�o"=菈Jj�����s;��-ÛX7���l��@�J���|�0��-���A����P�_�}.�ŴI�;S)�=�pn�\o��^�H
\�U�|���~aGm���B�%����X�)�o��H���9P�xf�M�/+����ݶ�S�SX����9
���诶�WQ�n�B4nA���=/���`�<�5�2#,�R�B��I�^�K:!O�Bw�2bZV�f�~BU���?"Z�l��wH!�N�&�׈q���" ӄ4gdI�����|��^+ ި��^T�)A����)ӛ��%�n
UO�'�å5h�h�Jؤ���p����2y�<�����E)s7m�g�i�n��k��§r'ť@�>�H�T�Ѫ���}vXұp�#�Z� HDEPA�ʣ<|���:��dA/٤����~���
9z[�6�$S�8�B
$N54�S�|�8�myA�~*lU�2~�ү�z	���P���c �p�ׄ4�f`\��#� .Ӕ�#��U���:�{O��t�1�ϲ������jχ�>�g��5��� ��x��C ޔ@.�=~^�\�"!�OԐ�ܠũI�b~��ʧ����P.r�tSx+Cl#�:��n_�$Q@�t²����I��2ը&~ϳ�rbHO�}"-`���¦4��v#���y,�r��X:�/H'a��d�w�ʉ����I�sUK١�Ϋ��}e��Z��q�������-�t^���DBc,�"�quC�b��[����R� ������+��P�.2��$@wI	'�.�֡'a�G;1z���ض�y������2�d�>b,J��R}�67FMâb���rX6��5�AM'�{��5f�� n*2gZIm
���UW�m
��Kƈ+4�C0��H�Fnq��ֹ�*,�c58$��������`Ε4��SԨz�q0�����_;��Lo	Ϣ���N�\��]�u�X�(��	�yevA��g�WՄ.9�L�����1M�}r\'0q���ky �S�0W��Y�;Ωb�2Zc��K����O��w��?��ȹ�:��!�&+
zV��熘%������1߶"�����`�g~��mid2m��<�)��_͖1�>o��d9���0e+�i\L��<�s�P\Ώ?L�ĥ�����"H*�~�N���j�;_	�S�-
+J��;~jY�e�w؇aL��r �qh}����k}\�ahj���"�/?e}�ށx�n�ܙw6�!���oD~m#�]��,8R�˃�ɥ�,hUa�zp>�'�X�\_��Vѓ��[r���[_����e�,�Á��g�:����(*1��7��,���SR֨:+�^&��\�͐w�����Z_W��-灩�7�-k��9�r�c�m�[Z� ��Usz����k���ɑ"|bZ�
���MS;0s�1t*
ȇ�$�ˉ�áW� �'jz�e%4e�*Kx�ct+Mf>V}[�5�'s�fa*� d�d<�����T��zr�Z��n�m�XE'����U|�8���<��������s�˙)`��Gl�1oC��"���:\q
ͪ�#%���{'!��� �]\��HV���߀~���Ձ�(0�m>��ϲ�@z;�QQnh\���(����~�?��U�./W�b����Ć�k�2����)��?��J%�f*X��rC�s��7V�����1z�z�c˭(8M��V������KU�q���_N���z� ����Y�4�|�k�(�F�i��MMZ���m�z�m]�`g�e�_ia�~���ˣx�����do�?"�ͪ\�B�ʍ
�Gf�`�E�`\	@�.�K����g��l�*W�����ÿ���{��i��aA�<��Z���=�ơ�fpnrS�eoJ�.J��W������N9�4�=�������r/�6���o�~��
��>,XS�d3*���ُL�!n,�('�\�ۤbA�ma�K�x���;�H`6�D?h��<���$���c�ֲ\(b�f�-j2\��c��xfx�H4�_�L�4ݡǸ��L����8�[H�m<&�ٜ��l�P��*����F���C½}z��j|N�����	��P��Y�Ht2m���5#�T =F\��W��K��q�RK���ͷ�&L�� r�J ��C�}P�y�" �Y\�f�2��hJ�,�ė#l�Y��A��A�(Я�uk�ب?5��d7U=�_|�J�BŸ��]Q��ߦH�uk�����F0~v�P7Y�Z�x:#�d�B	Lq'"T��T7�����xEh�D*}1���� K2�UY�a�/�������x�J�>/}-��}��u�������@xW0�'�s�l�l��M�$�F�B�DW��Ui�%E��":P���F���-
u��+�$�����ڍv4���=6�`V1�V�����9r��lv��j˥�)"����1x��ᔟ�䲴����͜��!s;�-6G_ᨾ�^�si+ⱡ*(��n�����u�"x�W��?M�e��7�qU��kBR�%\_���|��f3A���G{(|�ԊX������e9£Y|X���~#�I����U"�G�f������<�D4^?��I}��u~$��_��MB���z�~ w���k����JK���t�sLxt^QLE0O�7z�_���CnIM���&n1vܵfW��4;z8
#��m��cu�xżFo�%�m��5��{�cGt��0�D���8\җ���p�];��DM�̟9}Pp�Wl�L3�1d}��kN�v@q��vq菐v!����K���J����?Q�G~Fg|&���- *�o��*�ξk���{�0a���R'��OfO𼒄H����Ɯ{�`�
��9���wfè�Aѕ�����w���QW3z4�FÞ�/;�Й�	0��)_��al�����An�(�) Z���v����A���r.���qm��s�:���@j_h�=E�큆��BR��bCۊCM�[^t��!{�u54L!�01?ϭ�;����[�6�q�9b�����fz/�`�����xl��j�6YS�Q��3�N�)���5@x�S�ć�@Ϧ4�m\���~�Xد;�,�0�b0��n�C�� R�djQI���:��g�%A5rr�㦎��>�2D,�Rdmk�Ů�,W� ����-����3{�[$�/ɟ ���W��gxȌ�e��|���GHw6US){;2S"�rf�#RcF|{Q�6`�]�\V��b>1�i�'��!"z<�[j�N�d̏Rn������[��1�kx�u�c�Z��dJR2���oK�}��6L��+��uJ�6j��@�R����b���ޗԜ���d�	�d
�y����.ڙ����CcK�UًrL*e��A��śr�68��&0{�r��ґ&�L��
`�H�i�g1�Mt�	�0����ժ�&�_�����@
���'��-�-�%!��W��[ƩV4�P
.��l�Dq@վ3w���u�B�����-bU�;�N]���V#��vH�[ �N�]���Z�f� �wW{�8I+��V�w��a�z���v�o���d3�֓h����_y?����܂��2�:�x����;��I�\#��4�J[�]�tz%"3�m(�>�$b��{�%CɺT���"��b���a���Z�n�cK[S� �+��cX���]6���N����:0�i�Q���j�M���5}��i1�l~p�0�I�y���˦2�	��Tl����$�ƾ��2c�9�x�E�¬��|�9͸3��ԱVL��G�&��&�g��n�ꑗ�<(ZYˀi֛���~�rt9+u�:��ѻj��"y��O��]fI�
�~�_����I�^��ȥ|�7��D`�vm�$��v��J�mp�*�� �7��MK�V�.�-@�e�⁾:�T'�#���9"1�ڼe�)� с�O��U�~<c����X<E�O&��SځkxVGO��\S�m�"���E��x�OJ<� )ܫ�uuև�4��Y9�):F2���98�=s #8�9R� 50\��NV�m�p�"�J|;�`�I�~~�~ۄ|��{C%��5��5��r�������_�\h�g�$��RI��=�&n���v�6R�fVh��;���2�M1
��E�� ����	u#����Aq��Qr1�v�Rn�뒝���h��|�	�ڳW'�LA������Ubɦ�bA�Z Zh\�����۬�.�لK�/��w��6˖�b����ݷ{{Tv� �&Qf����1z���N�������y�ō�z��f�}sX����۟��>��8��6b�][T����G��-��X��gʭ>AǮ<�c"��z�-W����:�-ݰ�f��֧�_�H�h�GL9Zb�K��%v��<i�2���
��\�cI!�q��������j��[H���E�����;}0y&_����T�՛D��nD�n
������H3w
�Hgi���7�,��l_GdxeG�V�=r�t�o	�uk��3bQt+fZ�J#�A����JE𼸫TY�ϣ�%�V�E����V4�E��Vn�p-��rV�;oX��u$I,���X������zbRY>.V����ęW��6�
�x�}me�/���z�qW�d�=��`Cъ��C>��=&aN�?�o�v�2�bu�[�w��%�aU�8�áO�m�
�3�N����|_ں<����hI�h����P����(!�e�Z�A�-V��/��؆slr˘����Bѓ0$�`�ɲ�HV�C\{��'cy��':�kiq�'3T�Q!oBH���AT4RJ����e�1(�,��A�s(ט���]�wǜ׉i6J�A�~|�ž��X�ʖE%��=nKQն��ss��K�9O�nz�>g�u�*
vX'�*ͬ���e��W�j��r���Ԧ{���!��T/\�
��c�����]=ޓm����g\�Ӓ��%|��� `�i�5 �k�*
I�ǫE�ޙ��noAkU��c����<D�]b�w �K!��Z�Н��Ǿe]�!,h��_���\���/��>�rR1��Ii�3�g�Ū����pk@�D��Tw3 ��}L���tCC�l��p
�/�g)��"�U����͢��Xp�Z�t��W��=�j$Y�;+�Q���������Q>�A1:�y1R�յ�,���6��2���e.8��c��H&�Y�Ҋ���Ci���S]�7ί�Zr��K�N�AM��#�D����NW#��
�(�뛫�q����X7�B�}>����ۇ�C>����e��SAC,4��K�O�Q�ϊ��~U~B�����	,[��s]<�V i@�ĵ{�s��X��Q#!ȫ��Ln�M�bX=�7����r���G���d��R��l�K�$���0�]�|��ϩq�6���6Ŋ��."ċ� �<T"�j������f���v/��/�+����i��5�7�>��e�ktf7�����<�[P��I��֎v�͟3���nUĒ�~,�����9�~Oe���
�<��8%����E�P��F�-lϺ�)�E���['�Q8[�~���@��ћ�8+�'�'������mn~ƭs!��e���^^-DT�Ut�g�F�Rs��Z���?����!g�����%��r�D�n: ��E�c� zlߖ�t,�����ȯh�	d�qq�w�S���~J:���ߺ�0D�q�)��"�\b�I�G~�t��l�T�x2[_�0`V8�M�0�"�s#`9X'j_�Çj��6~V�5�o��RY5�k�I�<b��9�ԍ	i�����+	�&��t�e\�&u��ȚQ����i�C�%��u�b��ϰ��i�F�<P�J��H����@�G~>�+R�lJ��v|�����L?�Aۖ���4��_�c����,�Z`�Ө3�s��D�H�n��E�#�S���xT嚇���&����������Rzl_��	�y>}��f���,
��vZ�Gl�����B��YS�1�x�}:3W;}
�(o�R���*�å�+��Fm�ð��FD��n�D��K!pw�T8t�ԫ���Pb�ѰU?��G,��á/I��)a������ݓv�E��]��n�	&���|}�#yG�5���v\Td*�j1���F�iq�Z>Lӿ,�s�C�SW4�sB�z�����NPC�A	��!���� ^20��$Ϊ;C��\�>B��G��H��f[Bc+�Mi�?��̼x-��yt�C�ć���̺��f�ҿR�f-S�H�!�p��%�*���ｘ,��L�F?E�3�젶����Je�b�ֶc��銀H}^�g6qRƬ^s�h������� )�:����ۗ�d��\//��\6s����	�|��fժ��EvC�N����g�(ֆ�l�y���|��� 
�E��WF�����O���TK��պ��� �g�t��ѡ�),�Rt5%��!��![�l^�?�� ���'��OT�Fn:|�iI����nW	��$)堷uWV��l\,���:]ŨC=���H� �OkF�l���	�Ú�1�g}�����7��9����ԐN�*. 
���� Oݥ�}��N���5�C}�`�q���'�۠��J'C�<IՓ����4�w�ݜ�k�j�7c����;Mr� �6�����(��#= ��;����wɈ�	{�sV�O�=׉*�bV�(�F,�YW��:����l�Y:o�qFhf����q��˭#�-7^�9���GO�f�8Ȧ��(�����_zs�b��s��:��E�����7�Q}���q�t~$�(��?�Y��/G_��̥�1����Η��6㏀q��'F�B�`ʾ�U����Ø�&�����t�Z&��4Ӟ��=jeg��;Fʎ�ú:�Y��s�Ϫ��ܺ~9����D���
e�o�ֽ����L��2��9��%>�rN���mќ�S�?Vz��Y���M)Kn�^�P�>*�����l[����gTQ�ݪ�Iǿ��J��MG2�Z΁��t\�p��pB��8�0��j)������T]�;
��U]a�f܀ԋ���*�I6h-rj.���9�͘��V)f��_���`�Y7;�=�zw��_	+�����g��]��ƚ/wZ�.�[����y�P(CY���k*]�E��gB�j����R�t�G�90U�S����������ٸ�'�r0]'ט��'-Y���)aw�e�oBq]�W���&�,�֡ނ0��6q�ͼ����'gRsI�͎��z\��ڍ��eV�K�r2�q-c�x�7j�]�2����������?�_"�x
�ag�&);u�vQ�+�B)�����dv�eL���v]��Lj�O�ި�8���r��`R~FKr�_�4�a^�En��QH	�u�����U�}jy"0j~�r, ��/+y�m��\��nyГ��m#�-�y�c���]6鯑e&�Et���Q
^e9�P5[4p� a�1D��߅����˞��� �]W餹 *{Q�3D���ax�x��p�PK�0�u��7p̱	�[�O�����T�d`U=�R�'��Q�B�b���EE��5W�AA��h�$�oTۿ>�}lO�~���0�1p>e����D��-����}~�Y`�u�^�D�I�p,ke���|�:�K��ѯ��N-?�"u԰��DM��b����(>!�'|�y^�.Z����	UI�/�g��\�.
W� H����7���������ʤC��J�T��� ��L���>Y�r�y�Y7�v�FlQ�����8�Z��e,K5W���M�p,�i6r8�T�|8����2C o��a�>�|��>|f�f������v+{�O�dһ1�����,�7=� ��"����	J�
���J���(�`>��i�⹫�oM�������PHp���q��$c⏆��D�<)�o�3
 v�D�Ťw����`M���ȡմ�r�m��:~=�n~��G�����)&cwa5B\8�u��I#4 ���O�7p3��sC�0:�bQ�$���\���3���w*{8?G�u��`��n�y?��z6A�$�ez�K��Z;�'�2�W��Ni��7��5�z�����D���V�ط��6��py'�����7B�a�vs�M&_���@���$�s�|�XI�;�^�8��Բ c�)ɞl�4`3Yy��IoM�ԣUx��..P�*Əs��3�$�Q�*}�[_ToG�i�~v�c%?[n��ͽ�T������8&ZC����<u���ɗ���f����mOZ?�S�~�P��f���\<�����FD�Y��&!�h���c�I>o�k�y��Hv|r�(�����%��l$�iT!oh�`�A�6�d�A}[A��;<�m�z����� ୓���u���+	Z�r��Ӣ��ݛ��D���7��d~����	�Z����!�BPU�y�S�j���$~v�n�7 V�촽7YZ�W���eˏ�A?�%g��%�[}&�tr�c����YK|�u�c�J�%��S��m���� W��E��Q����@����5;1e^A�O�ɇ�f K9��$[�йe'���?���3�a�|��&��e6�}�B�4��sv�(���`��>s��Z�����	�����8����)�� ��'C%��nb-4Y��Ȣkˏ~��H�c�9��7�������Wg�i]QnfP�H���A�Z����wǴ�����5�D��}�� �Y�GF��:�b`1ԯ�v�B�$۽W��F���Q<�%��H��ή�_)��H{ĥ'�;��c��ֆImR�����'r'~�9 ���1�ҽQE�@ \}�� ��Y_S�����쌺�d�������1�_YI>>��Bb0M�T,:�o��S�Σ;
��ڤ�+�."��^��zCy�������%�h���8�f��aiѷ�Hm�����?�Թ����5�2��zl��f}kGl~p��l�+����_��y;0i�M�ܸ%�g��%���#�����_�H0�n�
q�yJȇ�4��l�� �����a�FO�˟Qp��Y�4�*AuG�NZ	��=\ ��J	����J���T}��)�X�P�7�fH+�����ܐ��3�����r�T�iC7���ʚ`)��D�z\L�4�o�'�ɉa�")Iq��VlV�6�f�D�JC�v;������{:D8�a�f�)���8��dk�\�lm"�@��D�������bNk,����x�N~���L��<��f]B�D�f�=��W�2d�[�{]ǎ��9aG/D��D��j�"<��\���p>��}Q��L_�؆ԏ|"��jG*��J�\��!V�*���z+B�O��Wv��A?AW�;ə�O�1��E���s	��NK{|�½�X�	��<6�O��I�W,7��~ys��4��_�Xۯ�#�Q��m�]����Ԉ�cp]ϏΙ�є��k,;��A��E<U���l���Fq=gB䬋�H�/Y
���1��ܗ����=	�LF����onHђ�rT4���P4����lh=��d����M�R~��T�̗j	�h���|���].�C��}ݺ�����ª�u݀G�Q���px]�&��\C���s��CƇ�s�K�H�쾪���z�S������.�X܅��Q	6�^`�����2���*�D���_�"@|���N�Þ�D���.�=�l>��A��?
n�h��v�#�~/��E�|���5�>�l�~��s���|B�e}$������y�����c"Nbv[JoJ�X�c�*}E����U�������M�F3��iB�����z7/�{H�����������Ν�������y#��l�wR
�[<���"Ϗ�u�:�}H����� ��A����E�r?T�{�h�J��ƪA=�R�\Db+�5suՊ0d�n����u��,�
�<L���͂t!�	=�v�*�	�	d����lX�S櫌�UR$�E��`;g
��O@R�$�)�#(lv�r�����:�H�7D��o�.�J���,hvg<&���>�o��\R7	h�l���رB��ДІ.+v!��^��^�� ҭu�5J�K�'ĈC�A}w�{�6��$Ԝ�]|\���VǼ�a�r�k�Ȁ��Ușs���ِ+&�2�������}��	��$���t��o�Gu�O$|�X�V�C��p04�{���<��0^"�]j����Խ���xm�pIz>r<�/`�!��a�|�'�-�Hux��s�U-D�����乿��I��ز���MYʑ]��؇��Z>�H!3:~�ֆU�� �C#����sE��i�p�CU���
�"���Ctw2�m�O@�x��Boɘ����X;��ŖF�1P�����J<�س��g��ݨ�l�Ͻ3!�Ċ��>?i�ʌz0s脪�:C�B;h�W�:�� ��<�$O$��D�q�	���¿c=K�=���X��8���ڼMv��-�*�὎x��3�2"u�Z�h����s�0�,mYh~��u���0�h�Ύyk��Q�]�x`]���e��F��� ����Uoށf\q0ˈ M`Sqzyw�,$[���h\���	2���Kٖ>i���L����'���}�@��t^{����Y��s1�]�vi'2�Ra];w��R���' E�W̢a=��R?�ܠ���>1�#��n��7�tx97�Gd|W�d�H�w�h�������o����(��ڈ��k�I4q��M�j!�X+ƅ���w���s6+��}��?9F�3I���;S�C��?t8�u�x���/N}�����yT[*��2����_s⟄z�7+���z�B��f���X�����(�RQ���G��~�&��<~>� ���	��^
A,�L=B
	�����K��z5��?�I������}ܰ<�p!%Xq.�U^���gh?��[x� x��D�Л���:>#���rX�zޖJR��6���j��̧�P��<z����{�{�O��6�����r�B��my��A�x�����iJe����Y	��ǕC��r:�x�Z�k��k�;ד�eEx�MrI������**�4�Q��K�-x�.��FZOYj���t���R�%у�W�Wb
��>��u�0����VU��7�K�T�������)�Ք���apZGbx(������V��,W����}&hy�m���G��4�s����b�A��`�~pe/�l������Y��ǣ'�|g��="��W�񅐟��h�9`��Ig��ok�a����2N
g�	�	<=�RZ	�1ەSӧ��!�u��FF�\�������*/z�9���#H�����)�2����rȋʴI!�,���ՒQ�x�W�۪�0�z��GT��˓pX��y��/5k�#h�=��9����S�'`6_0$7C.�ĮF�RZ��(���#���JK[�7�7�]��J���鯨�����k�8��Z�L�� Tp��!f���Ms�WXh���Y���+�>_UR]�� �{Ȣ"���Q���F!-I䒒!j���=0�v'��@�����6O�&N�F���L��/V�+��1���S*I�w}�ly
�C���--jz��g�R ~���[�qp��!^�U�9�\�y�ܳ:��J���oP;[������v��X���B�G�#��[�t/��|>q�qg�L��G���]l�=�ķt[g�!�g
��v�
S��;b
�Jr5����H*��Td����_C6���9P:-S�f:#gI��WP�Y}�qwGq�8/Q�qy�Ӵ�"2����j��E�Z��}�\��'j)j�Ք&�Z>�����T���?`�g/ ����#��(ɏS�Q��8���䙍N7
&�C���6��@����i�o�9�_�}Go �%�Q��z��_1c�/���Z���ϿbJ6�fe؁E�Ȣ�Sw�MTRu�}:��"�"���2 �+�C`�{�o�n���O�k�Ns�L%7��Fu�p|��0������~7�6��J�4�e@ �A�>�vs���������d�P^�K���8�0�W.B���]�(I�`��=��8E��6?�>�F*�O�p�+��T���ꄫ��m~a���0�h@Z����� ^������.*iT΋�/6YQfͯV�I5]�Q�Zn��JE�`l�n	��/���X6(�7�PҵކR ��p6�ٚ&���uT �<1r��,6?𝪥Mș����<�G 4Ì����-����;��x��#�o��t_K�+
 9��8�]Y�`f�-_�(oF�(�L6��Ā����;Zǰ[�k�"
�Un�~���̸�=�	�� �*��ݲT��<���9{�tj����4��2�<�޷3�� �g�`2vK>��~-���/^�Uq�Ӂ?_�W",��3�=I�����0G�����-o��s�ɐ6�x��Am����w���8��i�XG�͌�5�B���+�,ν�Vg�|ڱ3Kl�5t�_�o���W�PO՟@9T�:QH�@Gΰ;I2H�����#�{�yN��].��j�R-����!���1VR�I!|�X�j;x�xK�|���V6��>� )P�@YCh��G��]Yٮ���5݇+}����&��.��]5�?*�t��Z}�����m� *��j�f����`5aQ��C?�N�2�$�y�*����+����C�;�K-<y�*�aF���z��W̑��ڍ�K�Q~̤�9��&�W;��Ad���1c���i�jN���Ɣ��<��ܿC�}Jl��ao�R�%���6ǜ�'�ހbg�'�4�+��EQ�ڏtM��z%�1s��_���tZ�ht��*v���q:��[�	��ͫ�{�;`���Vx��-f�SP3����>X�!�ƧM�ɫ����C�@�9[J�Dw`�Q]o�o�HE��2~�cw�C}��ߪ]m�}�Ȅ�oo{v�W!~�IZ��}܀D'(�q���
�N�~@���������E�$ʀu/H�@���*�@�53�,k�0
�	�nLCQD$��XJ�>��L�p����u��cS~3�-�4UJNx���b<+��4��Mз�L��{�!�46n~���[] _>uB2���xX'�<`+���%<��=�^�K����w�ⳅʋy'�֕B�=��%E@�-��A@�7,��SU�����ml1��n��5O�T����,����ѷ+Пx���u�vm)��M$�|�'=�^�܀xJ�e$!��Ъ,�a�E)��:(�̹o����Ƀ�0[\�����#��d��#�qm��z[s���[�Y�LǾ��<7hX��q���b7����Y��3�:�7(K�dS��p��3�g]�U�,%�|�{�K'+�ЃAu�,
��J��)9�yU�i�>5�S�,m���i� [$���?p�\��,��^�h��j��,K@*���aź$�g���K�o���p��:�y�����'��F�vi	��xɏ<�	�M�v���4f0C%����k2 ���m��Ц���4
��ʷc��O����$��}S� �0��=
�MpG:Ĵ�h>~���h��>g��I���ux�~%"����jM���|ά��N��!�����z���@nʎg��s�~S<�zp�fz��8M0����o���t'6�X���g�g�������+h���85�-s�Pm�����N����,�����^'�m�|V����z��zl\�˽Q-��W��_T�?L�?��S	�Ѽ�E���aPAY��N�@I�S�nz�Z�b��ƖDt8��>���x�o�ɣ�%r%7.WW���:�:����E�m}?�̬��q�&c�&�!���9b`�8���r�X�4{{2e���0O�k��Q�ۂ�*?.�$#�APDJ�屗�[�W&�����]Vڑ��Z{�yԜuO��ݭ�g�v��~�_=G�`�ME�@*�}��Kf-ZF���9;���Pgߒv�q�e$���.6�V�0�芕���2�џ��NS?9I�kR-Fm)��d��@F}E��5@��d�DO���/��`q<,��j�YL�a�=�s�@��O(�lt�YD��Hc�6�)���R�fZ��U��^��1]�TkX9�����ZK�.��y��^?;V���~`NG������8+>H�������v.�q�{��Hl�.�@8��Af����G���~Kd�wꥮ8�
��Nے��_K� �kS��e�lkuv޶Ѽ��fzF�B]� ���m��ޏ�+�I���'(�<8>����d}vTL�t@<8�c�c�BT}mJqI�3��a���;ɛ�<Y�G�8p�B 9b�W"�y��x�^����~�|M5�Ue�o���)���q�������#�2���j7"+[��#��^�YZEN�ը@-��hg�e��m�F�������>_�v�
�(��I�Ь%`"]��r����Goŝıi<[K�3��e|
ˏg;�
��F;�JE�ފa�]����,�-w8m�P�=�r�h8�*���nu����4��(�M�ZZ�"�f�
*0��?���=��@^,�B��5t�>[.�[�sH�R�C5�J���-6>Gc��-Y�c��=�@9NR�xZ��AB�?,me[�ʪ|�/�k׬�	�_�\7�|����o���2OwichV$��+�E
�t+N8��~�i�
�2�f���{w>Zf�+��g~����WP<|��0���7g�bG�ֺh,����a1>(΃F,Ւ
5�`�8��'j���~$鍸�w��]�>��3ѳ8
`~MO4��,��G��;{�IU���L_9t���xh��+�:���`�?����n��ǪSv��Q7����N"��ڸdX��Mp�� O�lY61��j7�D�ǘF���|/c�8&X�|�!c�{Rz�Z1�i�|&`$���ߧK�6����y~W8B���\B`�dC _���~���Q��2"fn���@�sH���!F�հ@|d�'�Q��O��@I�O���J���
{ S^�s����иyn���
�X&���y�s�?VL>�BҞ�1)U6�~����k���]��~��P����mĲ�%k(�qGw�V\	��*e��Q��9r!XYw��@ƪ������(mt�١�q��Q�W#\�\����n��b��l�^_�9����\g�=#0��c�[ej�����Ӏ��vD�{��H��0��s�㲎���A��r/���ADA����>�_���=[�y)I��h�M[Z�w�����i�5
6��i����QJ��i��ɾ�^bC�]7Ԧ�ky/�������\���<?�N�Urh�,�7��e
)s��Ճ��5�����E��w�n�%K˨V�A@e����yz���;������h	kOeZ7}�86��>�b��y�&�K�����n��}aw�
���^9�b=��V���;e:�Hϱș�:;I�N�^�u�7�n盏Ӳ��/��n&H���^�p& ��&�G�B���)g�!p�X�jw4����LbqW��2J*ǝ��es�mׇD�=4���0j�2*���	4��Eί���W=E������ht|�ߨ�<ZGM�HC�WO��,ْ-v�*��H�۞^gE�K�v}诫رV��1�����#s4���;�����v��	a�m48�ɮfi� ��Y�j@67��.*UcVst�^���	�������uxs�Z���r�I�;��a3��dϙs�tiFM*���~�r �v}�V�
?�{�[�,�s�;p���J�8Ҥ�rePD��D?�"T4(CB
��[���~#
y|�_p��>�F�P�"����*H�5��Y��x#�a?���qS��D]m|kMl��엊$�~�r��w[5EѮsp
�s�>���'>�z���`=���E��%Q��N�u���/��"����`��ņ�^��?��P�rj�4��+|7V�)˙L�ز�J�Yk��x7/mHJ��+i�����o��T����p/������{O��T����u�]��`�|ޟ��HY-��;�Ԍ��5�II�@b�E_�C�+���FO٪�+�o�\���J5��`����*����,�s5Mu��5ӃU�Y7|���^�P������]�v���
����k7�*h����ٿM���۰�������\�筰]z&�i�j��p�x=���/.�qg�-g�'�JK���Pd��p7d$,��åȹ'�"q�zA!��p�a���ԸS��gw&A�x��ѿt���.�x����i1s����H��p.�,�d��M�tt�e7eZ��a������!M:c�.d[�}���5��Œ0K�e�2�����e6�'��������m�[5R�2Q�UAA-�qkbxp�t��K�Г��A�� 7�����L��R_0��c�^��(�R�#n�Ş�����=����E��P|�l�i}}Te��A��ev�/kP�ᑣ"Ғ�1@�=����CL�$tŜ8�ft��,�e�0T �s�濅�D�乄1C��o���LC����\rfJ@�S��2�K4�s&X�2�>���_(w{�=�O���<_�؛��`aU��cuG=g2��v;���p쬕a �ɍ�����[51��2�^���G��j>�
�z$u��+Th0|�"N�����6��dP���t�ۭ3��ɻ�p�wG��
P�SY`�f���s��:�`^ r�H賫6&�a� L!�VdJKN��dn�.(1�Z��4O}p:=�7��j�*8�ַ�$��2*`��l�|��2��b�*)������˰{7��aDg�1ʳׄK ��b� ����;R�ܳ�;�KU��A����H��E��nJ��o5�^+[9�(q)Z��<u�I�$����[�veD9䮵Ataش�[I��7	����O�dHl��#��@�+��Nr�u�#�cR�7hRAo��k����=�7q�Ttl�tvԶ�ӜK�G�J�@:K�"������T|c����M����_��s3���{NkHy��)Tԇܾe�췌��?;Np���L����L��;0�S��&�ejhu���=�j5�L�x�L'��Y�/��ZsK���J��w�m��,tXVR�M~ͳv�F��~��C�ͼ������B���T�50��Z�?c4$׶i(xM��~:(ݡ�Is���  ��n�v�j����il&�mCtO4�c�2��5;"��L�vu�L� d_T,<�`����a�~r{���"�eKe����!�~r�mOi ��v�g��B!4%����vb	�6<@E�ݿ�=!�C5s�+�*��T��%잷���i�T����~W�Cd����]Ps��q�$W�r�br��m�jY�]�a�b�S�2�UoXEe�����xϏ�4z2���ylo~��,exT��,�	O�0��!��?���r�r��ߒ���O(2�ʘ
Fr�l�3F_��Xd,@�T	���܉�ɧ�g�����.��W�g���ٗ<�'+'ZnӅ�/�P���H&ڕ�fx�o�JB�o�T�y@Z�����B��DmB���%�J(����ȫ� ���Bs��d�R���R�r�̬��-�G��s�<JKl`�,�4��=g��I��h)��"��
�,�}D���TD��([�3��|}Tx/d�X�� 7���u)�M̓=�`w�lV`�Y��6��;�Q9.�Sp��ᄣ$49S�DY��GwV�ͧ��Q�w�I ��]&1 eT3�^.��䃱����m����$�'퐰�*c�=V;ZK\�YjʦFx��au\%��N�]LvyU�/��W~�7j&����%���&��՞4��EA0�}b��,�PgU+�����yD��;ky���SS(6P}pv��e�b{�,�UӜM4*��:]�S{�Yq�z<�2�dq��w��{�~���2`�7���r�����AC/��r�8��Cc<ɘ�w������.P#�᫛uТ�.�-�������U'X&�M�H~��IF��	�X��(
t܆��yaet�A����kW�0�aCqԻ���Mɟ~���;��Z
�������v���O��¤~'e��09?y�qP0�' 8g�噧����Sçuw�)�Q��E�5�Bݩo�7�;;��$�EQ~+z�p��E�97�J�b�w�X�y���t�Ĝ����� tn36%�ec̔�b9�)w��|@&5YԵ{�bB����exg�N-��J��#��t�Ο�"bVE���}�G�/�6
6�ԖR-�����4�%��2�!��gȧyᙥd�����+��������$���~��#nW���08�C�j��{1�]�D�AxI\��JP�РTf���7 p�}�����vH&0]B��;p��hPX�J���NU���?��;H<gn��k��?�& �%{ ��N�\�����g�S�T���#,��/�w�&�D)OK�-��~��sA��,�Y
/�Έ�tu�S5��/
7�^�����5�}����V�a���u����_<��{�&�V���.��s��Ϟ\s��<�[��i�ʊ.}
%a�j�s�j�v~ܶ��׿͎O���ˣS�ti���b����X9}�vM��O���	�+���)�\ׄ��͹�P�P���+�8�V��+(��,1�4����f..�����e����@�\����W"��f"�!�'���#��Cq.�Ͼ��~3_��m�g2�������_��/Gn�]� g��(�I��.���Z�L�_�LH��;>aw�T[f���iI/�5�9�����pxm�����T%V��K��
��,�Jˡ�����p�R��8�#��	&�q�:�U�K
�:�/��Qt���k�:���W�V$)���Jg��ŃV�5������YZ�|�w�*e���O���U��T������zo��	�6�H���/��i��?��d�ܨq�([�r� Bہ!"�����c�sv��a�Eo{b'���fC�i�j�k3��ܖ�����$2�:a5��me����"�֤HI�rt	'ѣ��9�(^�0�=��VE@�� VuH�ՙ�9�Cs�`�Y� +�:T�#���l|�� ��p'�d¥x\�9�~_�~��u<�vSM�ܖk�����<���-,�d�٭{�nB�.��{��_��P��	E8���q��7	̟��Onqx�8�<����7�H0)�Jys���܃T�@���P��A
�4�����9����ʇ�q*�$����T��jΗb��'d�a�w^�Ih� ��g���k�k�ܖ%h������JY!��H�;)eaz��P��d�4��H�~sL�B�2����9^�C�I�l��]gA�P�<[�e,:���{��g����9z௴�Fڳ"���(	�=P��(3BJh��t��aS#1�� � P��^&G�6�+]�rwA��z1�5[��Ewv��T�R>٘�H�^��O��S��&�K�kIM��:�@r����`�~��6w����eQ��]U<7��u8�t����R�7Z���Y ae7Q�!J�����վh�����QI�m��o-2���¡h�5�{'SYI�nD���	�u�5C���9���at�\	f�!�e�3'���Qw+�[$Ϋ�%}�T�z[(q�Y�P�q�ut�tU��"����0;�_W�&��#7�D�����V/O%`�<]�X�.�m
�kK�I%�x`��K���;ML��ʿb��n殟��0/~k�u�x�_�%�H_�d�G���0HwƦfk��UՔ�P�t�#B��IEb��.OSmV�	0�-�#KK���\�X�z5ٵM}�sյ�D���/���<D����΀?�`G^f���ƍ�:���c�l�Y,0�lE��y_;<d;gq���o�
�[�4:�Lg�����������#������{܋�NpC��~��1��	����ɔT���aw���Ro�nu� J�/ޒ)�"Y@��fɻ�h loK�T=	I�Z ���0u!�E��9�{�cU�V��}�������Rq������$��,P�����v��b�U?
�p|�VLa�5Wp�	6_#7@��RuW˟3�
��aʂ\W���ޅ���#��׍V���U��k$�r!�3�ٚїk�:�� Y��R�	΁B:�*SH�i��I��&X�����cE�4k�:��۲C��en��Z�U"�sb�����Ҿ{G���*V�S�&���A�masں�o��z�[�6R���*
6�ZO�{-Z�c�;�>���=	���������#�N%���� +⌼��8���Y�Y=	�wkE9=��C\���쎘Vg�Y�l��l\�)�Kp�+Ў��k�?:Ѭ�o�Hű��ɱ.�k݈*����J $gm��D�c��;!��f�}u��;�"�-22�Y9��W�/:�� e��3�êaO�h���m�X.�(��,���Q��6�����=)�[�8��5��K�n^�!o��0�����kh]?+΂G`��9*iu���G�yNY��)�Y���)4��nQ�'|�N��J����r�!KB���K/�[�)����U��蝄�>=��1dƜ󮦚oO���`��Z�Ӱ~Z3CոWr���֗k	�9�3�5�ZC{�W�`����Ԇr�p�u�z�ޯ?u�;�p���/�"��2�SK8Y��px��ڐQ��v��l��S�I���^��,q<�ʫdZ��>��~E�ɍ�!�M3%��ײ�ud��,��� �}���S�~;q<_�Hd��]�����RaD)%���:�G`_����s{����$&�s��kY�oF/�<�.�<[eѰO��M�/�/ؖ=�}�*��^`N���de�_�?��*�cK# Ke�k�kP�������C��d��6��"t�N\���-n���f�HI�5{�al�����<U�K�hCy��/:���IVʧ�&�|T,����~<mR&�镤{�*f��R��]�3a�@(=��6�go�[��� �B����A�׸M�P��u3'���T:��ٶI�BNu��[���*����B`<ȭ$D�2�^�^Y ��#�����FT|�b�3T�'���:&�)1���S��ʼ�%!O�� e,�-Δ.x$7�c� �ps���{N�O��%��7�J��o�@�P6@<�*�`971[�%���r�|odlB��6K�h���2�_��X�?�3�ם^�/O�'��b�F~��	��?����X�J>c��@Ky2�~u
vfzG��o������|6�GR3k��:�l6�O���7�WGߚ`�����w%��I����%T�g>"�50�f�f��{�,��X��1)Z��v�D\�m5��ps�}���D��F&�n{13����r��G�}��v���K�{�Mõk(��#A�X��RIʛem���}�	
9\��!ꨑO*��	��Ç�G�uQ"5"�Y���j�p�Ѭ�/��{�_Ϳ��!P�db�X#C�4�چ�F0�	�~�C��6�����u��2��:��*-ߒW���������9kV�5�Qە̐q5����^��&�^Q�;����I\{9GE��t?�NK��;{�_Nm�\���\Ӽ�����s�Yt��v�_���{RZ��~�y?���t,x�vm�G^�s�����vLgw���
��>"���/B]�*΢��4T��ÜfCB���Tɲ�$�J��Q����#�6�z����Oɖ��Q�7�p�`橎��v��P���5���	J%��l��=YIC>��B�G�N���Hq��mZz�nfr��@,�l<�v�g&c�ΰ�#p�Tք
�bLrx�|�YIbph�ɞ$l�4s'�m���j>�1!�C�[���!u�֕� 9R��,4k������Ќๆi�x��Xe�ռ��7�NAx�ܵ<DP�0D<�7�I��(��9����i��A�%�n�P?�7���_����=_,'0�w�B���?�
^u�]ٚ�9X�u+���S������w���t��Í�xGOn@'��[�+���$R���[�	2*�㑪�!6=�琻�,8��n�1"�X��srt�EF�7xE�}U_7�jy���v����R���[��eo����4idA-U�/d5b�,R�F
ɩ=O�%����׈nm_E�W�I���!q�
;W@��U�pn�][����(ؒC�&S*�`�36��(�pۘ�E�>\�]��p�R5<8�x.dBq�p��?�7?�nx���N����)��(�"�p�����i�/[*_��[|��R8�q����?~��ȝ�c�N<�.@�\�c�Npb��
rЗFb�X�n)����{m,"��}_(g?���RU�Y|��8Z:Ah��׮���~���'zG�LҵL�������u�*��fno��"���^N�6�P�6d�#�l���
��0�>_��*z�XVa_�QD��e�W=3����Ցp']�6H�9vFC_�ӷn�i���WY��@Y���n�W��jMMS%���V�����>㺲-K�b�N��\��=A!�<�%DF��3
� 
n���,y���5/�]VMۿ[h̋~k�kğ_����:�ND�}%Z)�~�DC�%Y�P$�V��m$M)�Z��9OŋbgN����Jէ��{�7�,�ʄ��o2��b�)�n4̑����!�d��G��#C��h����E�a����H���@E��+x�m��Np���sw��rtFp3�=�D�ݍB�jǀ��4X$6f�9�2A�5��N�c&Γ�x�p#���p�tѶ�D�� �S�B�����>��J��DFI�W)N{�5��~5��]&���l��r�^�8Z�T�1y�?�7ꇃĕ�Kwlg~����\��Hl"���b��!��qB�_n�U�$�oH���fb�w���	#��	��H��g�U�E���#�PכQlK�����QO��h�8�|N#�ט�}�K�s;���R{W4��ND,Y����;���z(`G��|�ւ{�	ѻ������v񼒅�oe�Sv�T]�<%}�R[ݶ5 Y���~��4d�y��/C5��oh2\F���Ԏ+�Vd��,NWx���[�ga9�5���if�����Z<��������_}��.�'m�t�oQ�Z��5.Tv� �ƴ~�:��`_#b��Tj3�N��Z~'����u�������ڀ��� ����\HWp��{K��X٧��+;Zh3J(_� ��=�TO:\�QvDw>:�if֏6RW�G��H���VH�d�M'�LC.�������|����pd����Y��5�-Է3�(L5����&	����j�o�Ȱ��f�{T1���;��}�!�ӊ9��kUyܔ�񂒹-�0D�Q ���۩������.Ex�'R����EXX�i��,/�)(K�T��xp~� �"�^@f�!�(��Ch�C���G�3�J�<�C�̂Δ�H7Ư�?�as/���q.?1�51�GJBy;3�8�k����s7��R%a��E�n��SB���?�X��
����=b�̅�g����s���M��.�xSe���,��f�-4E�P$B�8�D%*��
�ZF	[[i��L��G�e�A��n	3R-�#�P��@����߇�7��n}.T�jka<Ϡ�(=;FّԘ��$���<��7���C.�����mm�bJ�x7����w�y�MM��_xgU����{i�48{I�հ��,a�Ҹ����&/���o����e�^U5���k����z�W�{x*�1��s�׭#����&���-������1C������Vp����N�8��R�{�X�l�n�$M���q?�DM��$��pAS�.�$OB`�?�� �p���.��֌k�A0tҸ�}9���^�"� �����8G���>���vP��mϺN+���c�Ht7����/�x�(7�U@��;ػ��䒎�Y����/*��Ƃ��Z���G�&��>���p4���e�x<�o9X(��߷p�c����m�%������o�I�p�מ�qk�U�Bʄ��4=2lG�E\Ѳ��1���p��Z�����Ȝt���}�Lƃ��Xؗ����LD����?��nM�6L�k�Q������]�i6R�A���+������D�w�W�U\�5�!���kr��U f�����l<�HE�ë�X�¾��x������E��N�@�[&j�v�v��u�����5�Wqt�+ ��R\�Ju�|��U(����R�Hށ�U�Ϣʓ5�����)�Z���!q�E��*�{�M��)1x�nU��OøA�VX��?�A�M�gpJ��m̸�
��\�K��l	4r��,Ƅ�P�F�)����H|b\��',�9E�^������K!��>�(���ܶ�����X�ǆ�)>R��0���у� ,'����n��t�	/l0������ĴH�����!�6 3ȿ��������sf�G}��p\��0����.�m|`
�çq��v�n*�#����{���qIL5��07ӄ�i��=�J��>R����7��P�C�.u�ğ������7��+��)��Dy�;�&���z�ڰ<�=#X{��xp�J��2�B�/�QV~w��m�]E��⢎���C�*���ߒ�ѺE�]H��#�*��q3'�n�uQ>t�/�|��a���I���˓�j�A� >e�&J ��'�B�ɊJ3���H[m�QF�/���<�Q��)f����R���̕v u�aB��diǊBJ�3�u^ư�&���řB��C�P�ϟ+���Է���
������<e�P���~@��R[ߍ�<'��ڵJ��[,�l�XP|iF��N�Vg��v\��]�ߎy�
v]'Q�Hi��NhUhZş-��Y��M��,���6�)̷�������e��"��y����P�W�H7;D�%z+���P�E�}>�FЮ[��G��uyF��H?.0�m�-]Z�Ýh�4�Phw���6Ϭ'8��w�ד��߾2$�㭜��ʺ2����o�s�0�E�PƦ/<*C7�#�W�&kȄ����OĎ*���
�����[@��W�r[a|�N�wT��Y�!Ɣ��5�[��d�vP� "3_'�yH�٦�ng	�V@LW�+�4��?�%�}UUv����:VF���4�3�w��H+� ���"L��f����['/L�֚��CG���H���H�J4�����z�I�B���t�;��	� �6�?1BF���^�t�R|��v���z����:���@��INc�
0J�9Pܞ������s�i�y�
���|j�+�j�l��e[7�&k�}��˼�m�����8I]4����Ӛ�Z	8]8�^;�$� ����I2����0�[��"���Gi�GoG�?��L}��KG'���|�C�������J¶�r�:0� I�S�e�k��$K�}O=��!�v�	����;ܝ�v���c����˹�H��k%D���5�	l��x�>�	������P[k�P+����X��\��=8�f�1~cå�s�DPy���\��Mj_%<�0�I3�4#Ы_!���� �����	egxn��L^w&H��H�^� ��{k�������p�K7��{B��[Ch�̽
v)Ӻ�a_��ʧ.�d��0U�~�|��,i;
Bi�LCT�?-�qd��f�E!�����
�b��*�_�i9��k���O:g;�b��RH:
�4C)l�0P��Q�4��?��x7}�.���<�Dѐ�M�=���) %��O��M�oR�h�2�.9��eO��J��� �ƺX^bŲ��g9�����6�;a�;�о���I��~���ͳ[b�H]�/�t+�E�4v�nSʏ�n86)y!�eg��f�%��8�֘q$ϻ�jh���J��m�h��׽y�Ku ��[?,F��U��1��Z7G�k�Q�C�?ڟ�om�vl�"d�[�����F��2xo�Ϡ�`w3��n�2d9qf�k���zT?�"�m�QLG�
\��빴aY��4+rQi��I#��X��QX��T�:�V-}�|�	�|�I��C:�� f<������p���k/03!��a�H�~�5���A�YTVB9��<�gR�H��G��L��.�n�kۙD����>��_a�fdַ����d+�C�r�v|ivIV�-P_B(O�����Ǹ+)I6�K�ezo	��u��B��g	<����5h�
�K`,
1��2UJNDޯ_����{^N~��xX�M�ۡ����,�U�v��G�L��� �Dlix��h��Z��HӃ�/(�^f�-xv��El�-E�+���}�� ��P#:�'2������m�i:8]\��y� vX"-�~��@fD�`���F��S�B%��'b;OU �Vh5.'���C�0��`,��j��,�#@�L*2�(�)�u1�}U.8N�����b�ѩi�<:.���J���ͅ�t^�6����J� ��)t���d�)���Ƕ�vT��� Y��Y-��>)�B-�'�YU%wLJ��a���t�2�7%Tmz�|�.�c �RT�.,?\�/i�?:l(r��|��Bkk�y�_���?+�v!�u�`P�x��-�?�8��]��c��9l���w�����u�o�1����ߟ�V^;�br"�3T���t�e拮�9�n�{��ګYk�Z�͈Re�w
���w���U�e�¾r\�:z�FK�g�LH��j�&��RD?U��F���'��G.���P���i[e8VC���� QE+Hl�<{�<��fq˴+���hK��x��Jy�AJ�2�r�>��fU��K���k��Q_�-�n,����.!�3_Q\x�0P��_5�y�A��C���]��ot��m��C`]��3=,�_sB�c�<C�bDk�2dL����@AۨKu$��x+�͞�w�٣|�a�?��`5��R�;ؿ�Iˋ�S7h��0:��ۏ�mh�n�kX�9b�Ȫ
A���J7po9W�y�؄�K}��x�Z��et����V�by~�P��;�ݰ�_Ƀ�Bn���<�vK���&�m۽c+B�7��q���!G�k�>���Ke3����`6��$�8"eW�M���#����S=%~�b�?X��2��$��{w+�{�?&�p�o����x�.;���޵�p۶���`�G���xpP��Hr8><s�e
�i�P�c�>�w�q�G�se��F����]Ó�����'$s�c�׵�:�n!��d(��p�x*�W��!؎�7%���휒trV����	�~)U�~<Qޞ��H�aϞ?�x�hl6�V
ec4n�x��Τ��DE��d�Ԁ�tk�$"�m��� ���4��Rq��B�m;ం�ěn ��A&�A�s����y�=☉a���1 a��w	���2���K�곡\\��Y2�2M�U���"~q#�5��	��n��=�°{��6�[�xc,n|�/��?`�t���**�繗v������>R(+un��n��M�j�4k*�h�v�ם��s]�a�[r$$/d*<�3�5]hX��;��@�����g�q�Q{��t�@2�-7�
�ŀ�5TF{�տ��C�&r����K����ki���L��C-�eݗp���^1�Ւ.`W�H��n�3�e�\V/�~y�Mk����O��2�.q9��q!g
�e^>gimV%��1�kN+�s-?� r��A�����-�9x	ث>���H/����K��Z�ї�>�o����ʰ��������K,Pk�0���}����2+I9誏�,/R�l��#�����)�w�͔��{o�Q�;F�:�ԉ)[2��i������jz�]O����64��Ef��`M6�y��� �����8�r�i��5_����	ł��7���6I�E�YpA5����G�" q\9�h�t�ѹ��wCf�D�Er��Wܹ��%t�$���#��_�]a˭�/�R��)�y�QU>�'����C� t�0Ȁg���4��fF9���X_	��;z�߻�L�8���X
z�4�a�D��	��d��m�Z�C����e�ā<2Q=�&r�%XM�����p%*�:�9K�����dj���� ���-	�f��.�f&ܦ'�o;��������1��oN+ �$X"�A�AT�(΀��*.ky !�X�K�;��_��k%-��"��b�6E��s�^��a�R�#��}|$ݨ��O�ɟ�x�mF�_��,�н�j��L@�.f"��{��)]
�H@FQ��-�H�$��^r����ڑHj�L�nR�{��)�wC���O�2��h��ey2�d�Y�Q�Rk��0Gea�<�$�Zm�g�>�YZV9�04{�K�fL�cN�؅Kid�������d8!�����8��TE�Tљ7�z�����R�X�ԟ��?�8�ye���o��R�y��g�q� ��H�_FX=������9p��d�'�`�6�����c-�ym����֫�	��,;@�"�D�z�qtÚ��������LƗ�+�6B�IWl���2*,���_0[(���T�%0o����\��.�'�Y'�Aޭz�ci˙�]����=x�����K�3 L]<����a��; w;�6)���]�QE��%�����ca
��H�Al��y�sJ���k1)��~��^`(�p;S�3�0���=����T\!!<��p��9jZ)K�����8ȯ���<���Ǥ�I#>d�+�~G�������,!rQ`^���eN�_�>�e��P��ξ6���ɚ/x��J�}J=PE��kӒX� �LK$�-W�d��Ѷg���l^QŸ-��{  ���N��^��[�M�m�Jc�����3*#w�:#�a�y>��s�<�h���x����N�C��^�aW$-u�ͨ�E��/���'���'�	�@���D����dohN�_��>�,Yʘ����H�ϥ�h�m]ݵ��0I-D�s@��5PQ����Gr�a����NGWu��� D�a ��nK[��/K�LT����є?�]]�� *��2O�#�m������f�דD'M@�m���1�6LO����W���M�m�Gd�kx��nF�(�V�l5��*�=����a�|R$�{���%�D����MNT@��(Ei'���ʁ���	ق�~3sm�Kʻu�糖=�}�И�qo$�e�m�WOr�r?�ma\�����~�S�r���I�Fv������,p��Iƕ��%u�݆�맼]pR������F*�I:\9�0����Y&܇�m�V�(�������HQ�C��,T��q��ы��[��_R*��e���q��Za���H�OP�R&A�^�����7�]Q�+� 1eJ@MD�y۹t'�Ox-UD�-��m���%�ؿtQ�8��^�7�7sF�O _Z���g2�*��ឥ��PXdS�%��Z�]��(�S�ni�L~*$d&�C�}������)	�
�H{2�n�3��0��É1;�q�� �(Yv��M�E���"4�����׶315V�sq��W�z5����u�N'��O��lڙKX1:CjXz�BOJC���8�Vx�3(B�$�㹲�D��Z�-�,��g�V��ԅ�eiT�ߞ&��l�Y=հH7^M��>zq��<�&�(�wA��9ìδ��9���5�ͦ@`4Kf��thA�et�A8^v�e<�.D�j�Ѥ�������5��<�z]ub�$E��k����*��37�ے��.,r���0�����[���"���Ft�����쏵������V�`�1H-��P�4�U�!���Si����O�np��W��m+<����E��V��Z��FƮu�����ݠ&fc@�f��w�}���!��+Ya�{H�#x�ܟ��7�,#��;��.)�4�_��w�(��"5�,�2��;aA�'Z��`�B��k�:�EZe�LV��������q�ᵹxT�>�Mx>��ͫf ��y@�'�]�����O�a�o����vl�@�_�2�E=}b�+��# R����L�n`k0u�.f4r��;�Ƿ�	 �c3-]%�`�},5��g��U����dsi��]��{����S�� c#�S��W�)h�W�-)�khۇ�i�����/���'�v��s�|�����iZȯ�D;��x^=m/�f��D����8�Z��J������]O�������O3�/ҋ��p��X�`�<9�fe��3�����	}D�O����^�"CE��Z޷=}���Z��nw(���&fɴ��4'%���mKA��8����+��� ~gX��&`J�^Hs55T�X�dg>�T��^��^��y�|TfRt&����d�S}�r=am++�9o��Nމ��r��<X�=����;EY�S$�~�&l�AbJ�H�I�kI[�[#Lt],�3p�W�/D���|>�Rn٬�H����Zs:
�Cd�m���X��kF4uoE���_�H���kT{��~!�ͼ*kN
�ƻ�"�H�P��>��m&{u<�r�N��XW�ж�N-�j�G�Lh�|��?Um��{��R���ώq�q�SY�0ԑ�[��eEz����51a�����Z6J�c�鞥3F]Tu5�q+8����vFp�57&�����ecM�|~Y� :t�Tf��+��<��.*�`e��d���d�{-<'��Q������t�ԅxW�r�Q}�U®������O@d���U$v�P�p��I͘:��$TY_{
������b�`_���֢px��j
{�S/��$ߑ��LY7W]������ai5��4�;�`�h XK�� IH뿢n>%e� ��涜�E0.�Y�A�V��Ee��3(?£��E�6֎��,�L�� �e}�����[��Ɵ�@����T-��oM灡�=w(��/}��`C���#㢌��J�پ���vI'��!Й�Ge�9�������Fzho��Y:m&�E�w	#av�PɕO��K��qt�)��Kk�4V	o.��\��3 :��@�T-YQ2�� <K��"��U��7�	4�S��<�m�^:Y�[�o�o���1%o��-�����u9���F�ݚpD��e�
e��;\z
,l�Ҡ�چj�!#�,���:�U��mT!LEܢ:�i�/T��4Q �!V=`,_4G��b�e��#Wٻ-,oVr+�/��	�_N�e!R����1`��� ��d���7Lg�d��_�����iK� )���=^^ₑ�Q(%�sVv�ZE�:�Nd����e�.K���X�b^�iW�4���[�A�%��"��4I��8Hr)��i����'�¿��;X�Q�"��e-1��nXe����a!���
骀{EnܮD�Y�m�����/C���}��G+�0˅A�Ġ�l<ؗf@��,z�P�p���)���u��Si��p�	�ta�5��*�?���12�K�<�p�xz�L!���a읫��5R�����r,�F���v=x�(�E6	oEUڒ���?EҴ7�N�2����ِo?�Y[�)no����C�W7�z�V&z�ZZ�:!�KNk�M}Fʌ�R��E0c���P����I|�A7�D��G�Ud8�����; 0�����O+�@Z�u@L,8t�GD~��NC�tۼ��&�Z�`(S���p9kg�D,~k%&�����[�ȑ~�����q���2��7T/�Eҷ�'�8h�*l�!����x�z<�4���y$�>P�a�2�Gk!��Vۀ
1�����{l��y#6�_/�MK�e�i���YHJc����� � �%�ē��z�������'Mu��M}CL��=
\�Z�{p��#���<w���'Y��+06�4�F�D�j�o����v�E��s�^�$:��90z�`g��@�Q�H���Ƿ`� �E�Vˍ!��ϥIi����وm��y����Mjs�Q����h���vr���I�y�2�N�z;�۵�[��i{8_�̑��{A}�F{�Yh��.�,��bCL��~�T�9&���3�N;H�.3��D$�r��.��M$
����y.A8�ó��Ż�u�#-��i�>gԁ��x�'I�x� �{�Bc[����+���$��Z�
z��a����"|�,؝������ڊ�7
�i妼��n��+�u*A���́��1��k�HcjI~��찞��.ޞ�H,�z�6�R�2qlJ���>�T;�ך��)و� I��?M�e5���aS�2��9F��vY,��| �b*O�!��H��?;�K������X��H����x�:�[S�)F�J�#�N���9Mo��%{�LJkQH)�(���Z�$�i���R�Q�D�;���M�y����#o�Uv������,�Z�3�-By�[q6Z�Er�V>�}9h7IɅ�t�z9p� K����B);����Udf���E)�� ��ꁾ�$���-��"{�WT���*ɀ��w����Q��8P�N��ؕ�+��w8rG �|c|ț[y�|��󥙬3�������$�s�1v~�F>OEw[G{�-߬g�}mꉺ.�_ދu�6�Ą��i<^7�~�$�i���|~���,���f7�W�c�"h�����М�W�53�r�rՄC7�#��j%gT�!)*2%���|w\=F.��ϰ4�8��j�f��4wˠ�#Cӈ�S�A�!�Znϻ�:���-���?X��O&MO��MÔ�ٟ>V&�EO�C��K9�/���6�A����L����� ��U�ݒ���zV!��"�2���X�i�qF���#�C&o	f����q�:[>��	_P漶�Lڬ�˂s'v���h��\+��o�ƔZi@��G���k���T�F�y�`�怫����B⃊��ϛ_#��Sb����?��h6��wm�����{�;+ZDpK̽c��A<� v�b����_B�x7��ԣ<h���2�]MO!����ޒ�б`���@i�`,�.��������А���8n`��.�9�.��#a�Z���5(#X�q]дW�e��;J0���~�n�G��f�^��}*9��TSI�m�f����0�	���v�����K'��>+#�c44�>Lm�����FN'HX���dB	�8i��&�ّ���X6~�t�5�J/��d��������J��ދ�J����/���#Y��7���͠Ʒ8�2�@�$��Ӟ��L:�\�p@���(�fʰ��$�m��	��z0*T��O�2�TE^��o����+���=��h�����ģe6��g�Q�_�h��ȰʟAs��Ǿ|�Եm��{� �E�n�=nc�%o��Ŧ����Q���Z��r����r|8��*��H�{X*i9�#����2�o�-����Mq���}׀(n㟤��������`A��T+}�n��X��<����j��Sq�}�݃+S��O|]�����Y+���Ϲ|ƈ�s��N�KߖA\Ȥ����=��F��~��L���Is��7��p �&ؾ7R�ih{���w����`3�C aO0�i�&��*<A�N�����=d�r���Z�=ˢvu��������KV������:@�^NK)}��-�zj5�zĄ�Ҹi��Xq$ot�޷�{S�DN�r�L��UF��$n��n	��t`���:j�&��� �X���S���;�W�+�Ԫ�����(��x�����b"*̹��m�{Pe�+�ȌLpI�n��=l�G󊽱����/�Bo����ʜ�T悧�z�޲�>�PʇW.Pf�V	����RMOx#����|4���m����H���}�ǭ)s������s�񚜂�bB�?E�^mYՊ$�C���ױ��$�pʠ��ݝ�V�I<��o��Cs�\�_߹.˙><'���ֵt
�H�Ǻ=�׾�X�y,<y�߸�D��g��#��EV�W�6��ɻ�7�*1N,܈ڙ ��A�Խ�]�3c��Z�����^'��D�5���|���)����`$��>�˴ �;�Ş��Q�Ç7#��X8%��`������-�]�e��[��+5 �7:S�S<j���	��� �E��j�ߦq����>�*��k�m)s�^���^�[s�b���pP�#���<�Bm��0d���g�|�V�`t2h�Lń��L�5�Ħ�3<$n��v�nm]¤q�f}-�c2pv?N(}aoX|�dh=c�����iǾ�d<B����g)!�-@xZ�w5�X��<m�x?��-�	�u��Ƴ*O�ݦF�̖�����HQ�4�S�T��x�7��zeH����,b�%�������9{���m_;�萖�9R��������F���0%��(�y���+Ёbޔ��P M� �8�8ZZ�*��~y��x-����?�DH.X�g�پ��Y�U��07��0���Ϟ�����\]c�Uʽ/�⩊LGq#Z��uxkKi��&L��?�I�E�C�ky? )n����bNi��r���c�X2�!��q�?�ll�O���e�����U'?� ��D�4IS|N�B�8��=k�[d�$z�p���9���Su����?T̫�
��,��a!a�Z�BnG�\�w���G�N��V��)�e�����j] ��!-�L�*�w41=�y�5sl��q�P�?���w�������d�8�·����pi������g���̶��@�4�R(z�6�6�"��
��y�<������H��Vqw�3x4A��w�ߨ��-�n~�8qU�",UڤϿK��u^.����#��
m�H�UI<��O�Z�����V���Ý�m���o]C�kP�EY�Xm}���z�%���/���p���1�i�H\����F�2��l�6�w��n��s�\å7���`C<��ːS�˺H6�f��=N�%�$�d�G��1I4��'W��ɔ����i�����5%>>�KGnA�۶�I©&)�/�X]�*���i���Qk'fXA� 8)8q�j�t�:Cf�r�IDpx԰B�P�>;0�*
�!�)�#�&���g�}+��!@S��םR�}���9�T�a?t�rW�(Y㇑)�K�ƪj�ҳ8�gT�1������Y�����>�:��g�?��6`����;K�%�cC��c�R�U�ӘܝL5i�����j�@.�ω0tG��GR���dRe��!@��ظ+��a�f�5�wh��Uk��0�i�:?ـG�a�VJ�r?㈶,� ��"��5���G���e�'~�]VU*̱��h5m��4��q{,�\�Sscj������B� 豕�aˉg�4����7� ��0�U�H��7܈�A��+����� �Ά%C4��O�w�Nhw� 1T�$����!M4uQ�����v'����N?��Ĥ#L�g�%��[�g)���R�r�~���LS}��F�!�@�I��z.�����XN�!?��`�t)�ԅY���[��"8V�hg�r^����O���E�]�V����H{�Đq�r%<�zz?�*����d���t���C���*
�\���<�3�p�^�1��y��M�~�(4�*�h�-o���N[K�t�ܤZs���u����)�ax�a��4_%EQ���s�9���'p�~�sm�1��%d��7�1r�������0kw�g�MM.�pgU��,8�2��Mwf!�V�4�=����r��@r��~:�W�=~C������:W^[hM�4Ӿ��b�y��$�F���.�4�+1'M֮J��ӕ1�KCh.�"�@}�Ї�Z� b@�*ȇ�Ԛ�+:�߲/"*�8�rKp�������n�6�<���ٱ{W����Y�?�ͶK��}ׅ��Ƿ��n��h��W+5ɠ�̗m��pEP��]v�D�8S��;�����MU�N��/��4�F�?Y��s���]o��!�gG���
��1�'� 0�������Ē�'�ON���6�;��1v((-�6I�r�i��؎�v��L�%	�eM��*��4��I���o�X�m�r������!0
Be�,<lB�}j��l^I�F��Ŧ�J�-C���c�A�̼�Es=�)��FJ�j�d�BYΗ��[:�M��EC �*��ӜB�q��x�n�hX���ť�\Ұ޻?"9�!��E��٪F�.�n�B�M:[<p���?|��3�z����_�\^N�ΐx�Q����h}E�v.��U�������;��̷�z��7�j�G��IVqql�Fz�l6���;?����=u$�{%�F,���1R�Y����\u~5�T�#"�b�9$����"H���}�h�Y����>�|��Я8��Ro�yh#Y���PQ��)�����2�����1F�����-�ŧEY2)�m�@H�(�2���J�q�SԾ����n��r�^�(=Gk�4�lfΝ���(�Ի�:�)	|�M���>�H��A���?�池ą��5+��(�UV�@j������A���L(�@��ь��z��D�I��)u��s��c����̧�0�*z�c��$�ߚ7��e8�q��#�e�{�a�ؽױ�E����Y��xE2���������h��.Q�]�����d
�<w�!DxAa���Jb՜�q ��&1j��cOp+o�6B���~���I%rD��\R��_��s*�՜��l��d�݄K�V�ة�W��7�{�4�C�1T�4�r����2g�OV�~��+�j.ұ��o���?��)����<W�_!�C�t�i�5Ґ���7������L"W�7-
\�o�m�q�n���:;�68����F=�[ Hڐ�ʗ�	wu�����]��Xh.,!�K�&f²tw����OJ�z�����������*�J��dۘ��B��r��y��h���BU����j��;��"!��ٱm_� �)ےh�KXFO��k�a`ܻ���~JR�HT�q	�7_���s%����ӂ�Q�����^��0w�ʞ]�A�q���ţ=dYJP��n/����-�6>�R�𸑓/�ƘM��C�j�I/ �8�	�J��ʵ�N|f;W�$�Е��ZZ�c*�-�'��Q�'U?����(4�qv:���f&�@��W.6��Ҋ����;u��Ɨ-#҅iIE���T�e�8?C�l(��foY��+uK)�0k���kH4��Xl��y�Mr�j�|���=����0��~1�q�����d;�7P������VKM�����0��۱� ���,��G��f��L��7�
s�L�J�z,�J���$_��(3�fH5����V�9�*-��2��y۱|�4�s��f}`!��h����"}��՜��In^�0G0P�}=q�db�׌���\�&���ۇ*9�M �L�^�n�3��R�d����V���Y5)x�إA�H��#Ú�ª�&$&2&5�02d|��jcF�-��jg/����J��?�Jޱ.e"ɦN�)S�9_s=9�����F�1�X���y\lE�� �CiH��n��2�҇��c��ZS$��
��{�0_1���� �q��s�?T�O	��̄S�ڙʩ���72���uw�uign؇])�qj甍�3��_�;�d��䖂�c�)2��y�H��S.�0�p
A����Z�O�}�I�9�D�)�L�žR0gv�҆Y2��*�|l�_d#5������+�D���"���Ț/��o9�=FVl�N�"��AI$�nY.}�ˁ^F[���?k��r�~�2��qV��~���s Y�+Fpƛ+n+ф����VH("�p>@E�� 8ƨ2'" #0�	��}��_�~?�)�i�@DX1���w��*�&��	���iX�H/��ϧ
x�fE�� Wy��!�˻����Z�,J�z��Rm��	���5L�Ϫi.��.�`�ҤP�C� E�//�/�]��H ��2����fUj��UC��HB�+� ��q�rئ X���eg�/=�(��0�q1��2�9^{�>���X�����a��>�_�
�v���[*p=����۲�P<�x��V�va��'am����*�$�l7��vrVOׄ	7w#÷��3�p+Ԛ�&�*ݓg��z(�M=Bq�p����*��E���)d��Ʊ����Y)��Pu(�$	\ �=h"6� 9�Z4�� ��W8m�����F[ς���&E�ز3�5�Ī�_�J�8��`�����#����|�B�=��)>�U�:��\��ML�Ɔf��� ��IL�P)L:B��?v���6��Ҙ0�"TI�Q�_�p*t[�	�8����@���4���$��HG9��YO����Z��Ϧ��C��鞜�~���!+�9����G}�J�N���8~t���6 ��YmL	̘��u2;�D���4�Ӷ������ܜ�`d7�,%(�5g�/���zDaf��^r����ƂĢ�EZv�e6Rg��IR��[ }K�"-�f�z��s����/�-Za�N�W(�}	E���5�&q�\�"(ޝ|�R��P� �1∊���{���z��ҁ91�?�c��f�TH!N�)R�nK'�+�36ӢE/n'3���$��B^*�����g5����e����WW|y�����g���Z�H�3Yt���N�U�	8���Le��+�S;�E{�L �"����_��_gj���-��MI+���yULtY��K��> #���?Qe���c #����[v�zm\��6,xyq�|Fo�ȓ��=M!��vBM����T$h���㦲q��p�b7zR�\����̠,�y�͍����g9�l�%�KZXo�s�4ˆ��	H�3����p��4"��6�\�7�x�h����D�=q��B	�Rs�[ހ�x���[��i��Vh��W��1}�:��Y����c��V>'��Df�^1�7P�o/C?9>u�;姧��|F��B"�Y���+{�w�G�������R&un�~G ��^�{s�i8������L���-�Sc��<�1�yv	�y{´V�m�r��#�Z]�bD��`+BK5���_�:#2{S��߆n���)���5F{X�;�ܟ�.��T�e�e�b�`�0�,`�=��km��íU�����/�,\��T���<<�c^{�[#l�d ���O�i�o�6I���5��ÀAQ�sD!f�F^^�:L��(ߐ>�Z»C�(���-H�d�x#&~KW���Xݶ#�K�3��Oo��][u�}݅�y�"�0l�<�pp���w�bY�.V�>�)���4>��p��+\��,!i6�������v���`%�΂\\ú,�� �-�A���%�ʓk˵	�Lj���gxRā�oM}��;��t ��ȼ��;ĒA,C�S\oçs(��B0�<��iKv��
���	@s�n�$�7��6%p�"zA�`/��ik8~�G����Fe<O�<W���짞��[=�7�V��f�/��U�]OU�&�f,j8�0�k�b��M��C=�<�Z֙����Z���=�ȥ�r�����bHq`w�2g=s���lq, ��3j�\$���6�H���^���h�u��o��Wۺo�P2���ދ<�l�F֮���p^P;�y_y ٷ��.��
=�� �]a���qzu^P�16��UywY�D4������z����4�1�s�t�+΂L�Yl���~�9�X0���[��®ЫU�Hk*bK���\ݗ��xo6E^^�aܒ�9
�!%�����W��3)Y��6SG*!�D���E!N��^���f9_&`��+�;�����7�G}�`����s��k*�N�Ӳ���츿�"�G��è�[��ήO���&�>rM�ϩ�,��ǗNț��7jBs�=�d�2���/�[�Jj>]�'��*�MV�N!>n AZ��@��ޭ^��PZ�����@d8���C����%���z�]�ſ�A�);�P0[��ɚ1�hU�oCӖrHNS:u^�%�xÁ�FJ�a�_��?�T*I�O���!��5�/��1��&p���g�n2�bZ�^-3��!6�!\BV�V��䒂��N�Z�0ч�M����V����U�I�b�w�E��Rb����V8@���χPgAq�E�7�wf��+��һ���QĔ���?�`���x��a�j��D.�&^c�gN�V�p</�������#~�.������G�S=�@����u�Gh:�v��tj�ӵ-�)��2_pCOo�\`���k$�C .B���}��0:� @g�W�����8P@O[GU{��m����J����J�k~��s R{�o�*M(�|
���B�ی�d</���8߫�1i����R��KrN~eN�ف �M0Ӻ��p����_��T��M�}8+hMBR�oŦ\����`�^�T"^dA��Sz�pU�d*�:�=����O��u����j(��n���LS���H����"�|�y.���+	K5R��g�Z���?U͠Y�B@���I4�/�crc��7/UW��S���՛
��Ǟ7`�݋�z�.Q(��Aߎ*���p�>�UYV͇�a"g�4�|һ�1e����v�|��3��~�|p�r���\>����8@���aY�gr>�e����E���U���ݬ�0R"�>� �Onz���-���!%D����o�����x> s�=ث"��褞��'K	�5|߆��s�kk��w(C֙�l�{�n����G$k��k�ۛ� �ѹY�{=�xZ�S�գ�������4�V:�0�J�4\H�V�,H�.ڲ ���V�F�|D|b �3#W�,9��=�vZ�s����4��F���L�S>�v���o�/VM�S��/u��.�Lͤ��/��C�1�ծ"�7b�~b���O���,�xiy[�n^���O���I�����+O���D�$w��y >X���<��������Qa�v�Zj���=��B)f�@4�w�����/����p�ܯ��� HkR�*�����=�[u�N��A���TZН�[ß�W��|�p�D�ν�z7X��(�$��:���-��ý�{�	SD�H���ͻ��nxț���g ��O�%�P���܎Cfzz����6�Ny�60G�䃸�lX^"B�܃m�'Ʊ���>�ց�-��܀*
D���M�u���P8�w��ͮ�����;/�.[�}['C�oq�B���&H�L�� $�����暰�rK���@\��:�H�J�X�*9}�b8j�?ڤ�>�q)�d�+�d�B����Y3����؉�~Q]	Z�$C�s�s~��A9�s
E����*wˍ�v���x���e8�{ɂ���l&4�ѱ���Ek��b@�<��y���uRG~0)^8��5P��QI�_��[��� TM�m|�rlӣ����ϟ�s�����Ǥt��~����<�6G1�����ɹXt�!��I�`�vg1TW#T�����sqy�v�٠��W,m��B��g�����W��D��u��i=!/�2Q�2��tPW;X1����#��q�4�#BG�M�� �����g3/ܘ�)y�1L�IX�Zn8�u�*^���ɱC&漙Gf|°�.Jm��5?:�s&'���K ݬ��%ǯ�+)q^a-�t'���YSW8\X���[�r>/G�+���!��E�ޮ:c.(pA��jz�����^n�0(�sY���Ȃ'�>X�h�Q�"	�1���QJjx�U�WnLH�;u�śUBq���xҿP@	t�Q$&���M�P���\p���G-ڸ������ڢ��� ��E&�ɑ�0A5���6���P�p�9��%��4ɘK�B��H���\�/~˚mA!	��z0�'K�Z�pGbMK�!l\��qO�З��Y�Zaw�	�2 ���EB�V#P��SBx_��L1��L�0����88I��졁�}�g?.�:η��
���ڐ~ں�� �4��E#�L`?�ɇ����.f�NnBm�����38l��EX�h��4�
%�� +��x����[_=�IW��|��PGi���IdC��Y�a):5��Э��6�z���g��j������m�x̢`d�T?�hV�*rϬ�lK��~M%Nb�ƴ�7e���$��,�[r5,��~|kY�]π��23N�[�5F����w�K9�%ʆpn��g����X��ʻ7�ധ��srɸ}�9���,��NK����J��ES��~+���.�9xY�F���S�{@2oi�|�g)H
3���Va�R�
���m�F��G�i��r�m�AoF�D��bHH��E�YW&�� �O	��=���v�5������m;C�u�T����< �7��v��o8EY=��c	vv1�"{���`UeI���Vzh�z��N�so�����������r��S����z3Y�LJ�]�YԂ��Ĉ��9)�*�-_t*�?���H�OU��C��/Ȥ��2�[�o��Sd��_}�����e�#k@,2����Q)�뒺oU"��c/A�=���Hߙ���EΠ]�֗*ɱ����ݑ�W����6yPT���s˾"܊��7и��FΙ��E�|7ʞ?*���ǈ��/�cE�n_���<(����C���bP2ӹ.�Y*�8�(h�-R[7�Ѽ%h,Ylɀ���ލ/Go�� _X�*�y��p���N.ߞ"h�]R�T�(����@+��̍�M4�)H��^�m�W� ��if�M Ine�U��N��.+	 �����җ̹e����Ѕл�O�ڶ��ٷ�^k�z?~X>]�/�O[���N��L��a*	V	�M��z~�Z��|^}����K�Ĳ�Wي�z&f��zN�y-�TߟUn�:����tv�&s�y�|f��3
=Ok�����H��@3Q���_n_�1�
]��.M�p�ۉ�@H�Ѵ����ay��-�΃�J��i�L�B������|`�MB�̉4#B�|"�]�-A��
Ln�|agy�"�"B�xD@��!��YS�3�(�[y'e���l93�[�)\}'LvC��.��z��"�>�u����o�{�ل���;���`S���f���+BZ��K�R3|8��W���=tDx�Dlʋ`L�MU�(ˡ -�H�8B7{ϹY�\�� :o%��mFl>�%u���Nj������/u��T�P����Ӑ��s�M	>���U�ј�3���魲��I�)O|�ِ*��&b��唩Y�<S�tK��@��1i4Rf~b�L�`���rs��;�?��37�T�|�,�:і�MVa*�e\u�ᅭ 
��l;�XōF�40=�E3ٔ(�{
�$�;�Y/��{�y!�M���^"�j~�4���l�:����	�Er�1|w^���t��+���Tg �Q��H�'�6�#����~�:���H�	�rT3n��������r��H)�@�_���<T�F�ꁜX�}��8̉{j8��ٸ�<w�������x��9��#�#xlW-h�\Y�%3�	PlB7bu�v��Z�C���/@�!{�G�+��X���Z��pI�ny�%7/��V�b���c�(��2dY�p.��}�i(����5���EgbYX�󢑧J��4�=��yU0����z����/a˻3��kԐdO"�1G����Z�}�ܚ�A趨M��a� S��q`�_�r{D�:	d[��o!Y�g� dI�$��.g�wn~ws�/K60Z�C_{yw��ܚc ���5e����r�b�~������l_�B:Rt�,S���4�0h��`�F����$J�ǁo�m�AP��
�Su�KH,q���x@�R���'�{�i���'���7 �����N�:�2�T!Y-�j�9J%��������O�(�Rd����R'6C�i&8�9�n�� 1'�ďW�`»�G5_���A������ r���^��R�i����kS/&�(���ɴ�)�pWc	�>!�wMCQ�tK��,4.iU/],Q��(L�^�����@���V��.~����Qҫ� O'%��xSCk� �.w�!��@�vT��8/��qm�������|�8�+�ے�">S	&�����-˻�y��!�[q�"%�����c�;WF�3y�-/u qk�w[[��[�b�<lɦH^��\�}�W��P�ܪ�ԙ)�N�^��(.�6��E��)$'���M*A��9T�6j��G�Pٸ��K�m���"ܔWwZ�rIO��쥩�(�t�hSN~�~�_xO��N��n���5����7�ۗ�G�uݾXKW�@�g�')�3�wZa��S�@����1���J�'Jc�ۖ��>_ǌ2f�f��J|�'�]r������o��( �������n��bp(V�v����g�n.46t� �����*�\��~^�Ѷ0��&����P�_w�4�������m�|1���X����	�o�:�7D���c}d�.3У,���"��8�����b3�+n] .���Ď�Oo'��T��M ��D~W� ܗ%T_u�"F�T��3�e�c���׃f!$�]K��#�:ߒVE�r�uB�+��K� ���$��:�����L#˹�.=�[)���PCj���u=�|q�%�w�:��I�ԃ3˒��I�wR+���G�C�;���󻪫¤e�Pw��齀�Z�Tr~1
�0�����sJ���Q�y��nf��	�?T�:5U9�^�kEJ}�\	��P�� �. ŧ^�ta�X���qf%��"�TlZ47`�K,���ĳ�1�#�]�!Fa�KIܷ��-˛�M'�m��Φ��E�P3�.*�r�R�}�!LA�AT��X�B�o~�:���$�&��f����̞d69}�v����$I��������!�uu�ϑP.V�=<�y!B���F���6�>/��`���=����R���I�~J�@��xk����w�L�o�����$5tˈ&jx����4�P���N�Bh|֔�A�(�t�������*T�LI�)E�k�9H��)�M��m1>I*� N��n��\P%�H�"��P�fK��|���4�=T�]*>:�ҷ��ۇ�_���mqř��>�D��'~��/6�_��_��p��]lD��Ů��r����h���ҕ��	�����\�r�l���7S���"��wq�l�
�T����eg��	���'O�����7��VZ:_A�p~%u
\��: s�㍞:�/`��	�� �q�o���v��]��^'��A*[��ޅ���~ʎ{c81vUѨބ�?����@���1�o*�M;rw���u��e�e优g����%Bv+���<�˞�S`�B�km�|��.ێ�`���1ѡ�IVq�=��=Z4�'�L�Ե��6O(^��.���xY� �SvYlU�M��L���e�Lw�v���i�ftѢ{���)����`��!x�~;Ylۆ�)i�-�>�J��f<���K��� R �D08����> ��)�
���ս�̦�g|��YUw���<` �s�>�o,܉�����kjq	�ro��&A�x���}�D�k�n�#(�>MK~\� ��l�Ǡ��~<j�k��Q���/u��Y�����v�;	�N3��M�t�ҭ�qd8%�J�-��>���v���\��Q�о�,�� M�L9��#g��gOZ�ٕ$�P mT�-T�Y=��U��a������+ԊR#�kA���|�-[ے��rQ_p��l'&��L�bOt�>ƿ{��Ў��?�I�7�d�XX�2�
�.OkoYc`�>�oG��L�#�z��L?т�)�~�����ѻm�'�W�?�R�߉.�uy��z崻��2��>�Q9�Ԍ� 0���l_�FT�M���
�k��;��9[��>vx=wO�p{?]�R@oǸ��Ϛ�k!�>�{pBX�2�R����/r��GU�,qg7������mj
_�Q��e���wVIY)u��2ΔN�C�-6�W�p|�9��9Hz��~�zl��ikn�?��J�}ϧ@������^
[�@d�F��ZѠ�߯�߸r����@�4���
�=1�UI�����W	���gk٘P<�#����ѺL�Ʌ�1����D�&�����%&Sz�J|�VG�(>/�X	X`H�1F�?���7�t�J6��l�%s}w�Q���C�y�\N���*ob0�O�K	����_�(k�-0��s��K0���Gk�*�� Ce��t��0�-��OH|.���8{��n��/mЭ�=��UE]�{����{����]����*`w/HaZ$���+;��.��46���Q&����)U������rptUtp���}3�2i0���vj���I_7���=]{����<,� U�P��׀H�>_��d�|hm��Q� .��@�`Y�"`�? �}=�:~� m�4�3��o�髪-yoY�L��m�r��j��[���+�,Q':ܡ���/؅��8*���uM*�ő����?3~%c�Z.�*&3W���V'F��	Q����ˎ[�#�Jі5=��3�)^���|��/�aU��]����S��n8G��Hc���Omq��WRW$!	�RT��z[�ȏ�;��Z��h>�w�<�&�#���`>\ ϑ�IKް�sF�زi��C�۵l�XϷ�0�L�I��?��.
#o[x���Nt�q�1��V�.sU~ު�m`mS������n͸NܦW�0�s3�X)`<V@
l`O�?���ߎ�=�`%]��,��D�"
�qLj�|D1fD�V�Ц���db�q���!�NveW�-[�H���˭E
Rt�R���ݍ�L
�U��͝�t����&�pK���x�^�f@|r�,����L{W��5+���_G�ȯ�X�����E�h�|�O/2*�ϸnXad��uIJ�����T���4"B?Ŷ\EQ>��J���[ò:���8�4�{J���m[��=�"z�����dy�&�2�£pd��X,Z��qm��3ٷSr7?�z}K������T�Ű�~���G��HYդ��:o��r���C��,o<�m��o����Q��AKs�bO�����޸����%{ɯ4��vU���L_w�F���\~�<�i|� c�x���e��I�h*o����˛��;�)��R���2!Wx�(�<]o���L�0��mIl���X��*R�6�co�H*�$��G�̅,��^�0J�+]I�_�8X!�ЎU�<x��VT��@�Ш3 �s����&Wa��x��F��c:T�'�k\�Y|�
*�n��O��������n������`^x�<�|��P���i��"A#s�5��$Fh������p��Se�Z���d��NP�l�ϕ�P����μ�2g��2
5�.�r�#��8� �؄�z��2����_3K����E�[3:��'�ũ.�)� ���/[�P
�e0�|�/�5�7�Q��B	/h�%R���c����g�h�{�g�|	_��;���l_:ښ�p��k��1]>��*׆�)�Ā$��VO�7�A�{n��Ĳ�i�D�̼��x �b߮����:;~�5yH��i���H�ڌY���D���j#�x&���q�*W6q����X&_��Kܼ8j�r��$WŹw���ZG�,�G!�h�>� ����<��į��Ȱx"��u���I��Q=ti1~�؎Ѥ���$�+�k��D��#��V�:���g���"�"#�ɨ4df��(��*���)�ˈ$i� ��,�5�x�%�cM�ѧ��[�[)�Z�s��Sr�8��_T���ؼ
������l�e���^l���p��
,��O!Ssِ%�!Ϲ�.�`;�|Q��˯���Ԛ��I`J�g�Y�i)W�̠XKu����*$=����=�}����b\5woÎ=p��t�&Ő�X��+���T�.�j����s61!��Gj�C�=roKZ2� G�=[�ٻ��8���Ne���"�߹i�˶�S��僡j��H�;��+F�;�&�i���"/��_��!X�_m�0H]U�<3{I�=&dZ��O&/^�D�~����Ag�~���}���"��".q�'T���f?�������
l����+��*�lvE&��7\������z&��ٯ:����$��̜��q[Ls��uc��@7qloQ�N>��%�Y���K~�ju���-xu�TIY����~t�Ӗzϊ�(��1���;���_�ŊA��#��+��l��"�%��u���8IGk����x3�jMl��m���;=��Q����c�w�Mpc���l�_}�]��޻��y{��H�U��֐:���u�5n�i�P�vV�X�`�h�Z!/��ҙ=\D=$�.k��+����vst�0�t֫ )����$d�ql����L(�Pfk�B$̞3���t�
�]?f�=>\{}����&Z�n7 �����>$/E����R+�`����-�W����s^�r�~���V���Lv�v����^R�Cw� -�~��	F7c~3���s$S�����G~4���
����Z�6���!�G�}8 tucU^�!�j/���U���{��#���r�g)u\��A��Y�C�U��Q� ���~�����{��`!f�/أ4F�/듶l�^G��@�O�|��D���^����kL���=�n!��؄wj~y�M0��n
ɎZ��7)���c|���㏌mB2����a����+��'=�|,7��zf~��8LFU�g����r.�e��� ��kyOXj|%�Tw��B^\_L<����2]��x�$��҈w�҃6�Ҿ����N�������}�kA�,�-xN�V|�|W��;G���>F�t:�ߎ�/�8��p��)*l�FW�DtO���U�0/*���qc�V�!���B�D�J8�=��2KTCP�)�O�C������@�C����l��ޛg��Ip5F{c�~36dU�����7��3��d(�T���	pZ��<�q�k�sMQnG�;i|E>㶟��� ���4{]�U�L������^��;ۯ0��L&V��ZV��S*�+խ���- �۔�a_�T�m�t��qh5ms��G�����[�_���9t������P;i0�a�X��4e�^XKB��5�?���l�"c��՝��K�3����ŞK��|���bOL�T�˨2.]�e`5�[_@�tuT4�n�RX�h 2*5��gc��׊A��I�I�����p-���WT0�+�2���X������q�`�a[ގ��� ��~h���=L�r'N�$D��X�y�v��
{c��� ��}���D����lz�f�:���h�(d1��緞d\�<�yI���N6��9��W��D$F�7�1ͽ�D�X�f��X逸!i�,�ZB�BL�w��� cچ����
�d9����'d���P'�"}���pQzC���	9��c��z{��0hγ�}��=m�+,j�:�Yk��������g��H{�7�����d��WF��R�+i��ߧ�: :1>�LC���޿��+���kN����˵ Y<�!s	Go>�"M8k�L�.�^� k�	�ء�A��w�t�'���82AN`"P��Wi�M2�K�Z���扢{Y�b]��U��٩�x�c�y�(���i�%�TI�%�&Q�E����N�+;_��5�#��eO��x��$Ȅ1i�O'�T�(���x�)��r�fB��fjԈ�Z�R{8��J
A�	|�(8�9:�xʔ�C�jL�9���xV�F/+`��5<�7G�\��^��@5>�v�I
�A�N�3�;�%����a�?>rX�]��9�<g �!���s��a��{T;�[��w�Z�k� ?��>T�E�b�b�'�#�s!}y�U��?@�]���\H�4I�e��4F[UZVŔ+B�k�N؎X���*Ը~�"Y�A(��E�W�`���;�����Ob�= �j�����2t������<跳�>c�	*?i4c>�]�����W�����@ty��%����ו̉�NS`�_���K3K�n3y�G�R$9�{1�X%�V*
��9ң'�3�x	�:+=���C�)嘅y�<�s��\�gU�]�<)y����JY�sɩ��/�5C�{K�tJ0�R���N0�я�Z�u���TH_�3K�I\�@��!��se4�$\�p��ۭ_����q+��:��W���^*��Ѽ'���~�}����|w��n���D�qcO����NL�#9Lf)n�}�T㐋R�05��8�R�#q���X��Խ!I��#���H�a.�l1ʩw'
W/I{�e,BZnl�,D+y�ռ&ɚ2}43��-��9��p PQ*� �N`7��΄�Q���L�����Z�"�7]~LB�Z��N���js�xNC �qߎ~;�4�ɮ�/�rm%���o�A^�GI��q�A�:%����'Ɏ!��I�g�ܚSb��}�~�%����_�J�
x#CFUj���gjo�|�J;Hߒ&m�y�@Pqyy��Aa2���%l����5�S?�|O�lլ
0����.٩�=N�� �������D�mpR8}��S�Q8{L�����оL`��4°�qw@���1�#$��%v�J�"��u[�����?E�*��tj�S3� �NvLa�X�d[�%h���7���,Ĉ�Z0Ĩ�8�p�}:��\�W`�c���\����k?.�����ё����f��Z	`"9�;5�B`-*i��G/��Ѻl欇q爈jő^��:�vYw���#���Fx��,,h�s���b#�h����P,��l�s�E���<�P
�'�q��N���[�O4����s@b��s�N�H�Gʔ����rD��r/j3�!�~m@��m�7s�'`ɶ:FW<��D���V15_�}���H�tM4�ƙ��7D���aW�As��}j�u�[/�1���4II޵fAfPi��e4�=u)@��ͨ�0��'D���]�#>ǂLO�w��y�$���/7�Б9f{��:�J�2���*x֊/;�WZ�DY#�n�ĭ
+���J����m�oVӪ��t��f��n��
vK�P�W���w��(�(G���"bR�D���8ie(T��S����u�|z�A��Bϱ���;/s�:��!G��a�IC���t�j�r�-*Eۓ�����d��loXaL�+2 J�d!����(�?</ �Ή�Eb��������9��e��f�%�*�e�v�"ŝ�V�������5���1�� �:�:�~�˟�U��N_�FE�`��3M���k��r�@*�@%��M0�fǝm���Vo@_R&%��SkF���)���~�v�-����fmH:�h�w�<w2���n%)�ݸ��Vm�;���E�$Y�����y� w�PP�*��A�Qю�@I#�^�:��o�mϏ���ű�5V+�-x�u��7���"{��bP˱��n{�P�CS��*����;CN{�Y"l�Z�~��?D� Y��$��[�k+C0-�lЪ�	JwU#�_����["k��5,ӶCg[����͢<L4�i�����D�[���+�zIߍ�@Y����>��?i����������G��y������gr<(��n�?jΣ���|�۳�ĭ�(	����{���b���@�T��m.I�+�S(��L+�"���q���"�l����;`M%ʰe������׻ٺ�p�]�m�(��sS<R���*����)diCtE^��s�i+���-;2��
�-�����嶄�����M�����2Di�̴�϶N�ѧ���}�5`��m���>l�5��D�o7X׺Ԕ�����V�+j6�-V���!�7��1=X��W3Qx.�%'0pg\w&�.0ڮ-���V"�0�6���R���E��z^gs�E_t�f������>��k ��/<�)�{�Y��%g7w8�JD��z�=-���A��TS���
��ƹ�6��g��i݉AXF�� �.-��D�ߙˋXP�fr�Yh�e�M
T����j�ժ� ��sV��qYi1B��s��S8�} ���o�J�mǎ#��t�Q�I�l��q͉�'RQ�c�֬���NQ�p���A��z�~[�]	Ox�a֣Y�Xpq�
�M<�O����e�+�[���~ǭˇ�nb#53�)��	ra�e�j�p7�cǟ6^�i`.A�QI��b�t�8�-�;״Fa]ȡ�Ą>fQ�=j�}Ge�٧O�dV�Z=M������'ɦ4M�
VIk���g�V�(!��30`S[zDK��b=uL0j���:��>h]�E�ue�pp��,�'�l(�?���nw��4ۨ�&˓�qm;;jr&�'.�������/�;�	92��H���0\6zʛ8�k��}p�ǔe�Oԉ��^��NF�2 �H����zƑ	ރ���c�*��s<�=P�j��<�����4uE~ 4��Lbq�����꩘��0���Y��s� �g���������~xa'�M|����� �nK��E��?�����XT�K2�ƻK�i���D���x�>oÞ�������y��zk�r|���#Pj�!��.ɥ���[��NNo��Mt����{�2��E����gPKM��_⚶��xo��ȗ1���vw�����0��s�C�[���Ul�D�AR'��w����
T�2r��tt��B�u�*B��>I:Kn�_)A��+��0�	@�o�9,����.��9��o��I�L�V_�����8C���k�s�G�������
�����"�~>%�p�%EEY��;\�ɾP�Û%��j|���{O"����W��A��/����!S�����`��u�C����`X�_7[�&�K��D�W��ζ����Aʢm�����(��-�8L4���P��f�=�w�.1����7���־;������|E�+�)����كK�̝���`h�3!�LD������^̩FN�x�hF�t!���	0 '�c����~Dt�Y'-84�XM�:�c��t��`x�$7�8߃�^�Ƌ���MGϹ�ƮU:�.�$?CIy���x 1K䙮!w�:��"�X���uia�J8|)�l�����HG�Mψ����j?2۾��BP��eԕ��Qs��ԡX>t��_�؜!:�j[��vLX��[�_O��$���9�yG�v�,V5�w�S�[vR�(��e>�A�F���ӟ���E�6�3�$��aO��b�P�|�&�����s/�=��u��{�3��"CT����]Z�k?N�Q��.�63!q��a(�}-4����g�&��7�.�L�ۿ���gd�bC���cN�^ji�<�A���(����l<�4�&��B����m�N| �����.��>��Cd�z�Q��z=�̨�̼Zq*���v|wY876O�Y*)�R�z��,���@�׈�l���o�c̏<d�&�Q�sf�,��
�'bhZ�4�_9��̌����������M�`��Z��̄L�rǮ��qIq���II��t�:��L)DӺc���5���|�D�QW{�""@�m��-%뮸����W�J��v���j/�m�E%[�Vt�ʓ���f�[z������yM"��)zm��P���Y}Mɞ�����?��Lod���L���_�)����{sP2�yK��;���+@	��c,�sמtk&��f(t��ݣ-��1H����o�1���Y`uw79 ~c�D��׈�������6�f���GΖ�K-�-k[N���-���(���}b)C
u��qkS\���S�;���
�����خpGJ�`��+��y�>�8��IЁi�	�7f��r?���L�*�����b�B�`�stѸ�mJ�����q���H=X2�C#�� ���!��O�Ti�^>e\A�0�!�LXz��YL����κ�C�Z�Pa� �7^+�Gv�@�W�&0�l5w�Uͷ0n�qG��_ˬO��&���i�y<��a�f&y���~�T�H�b���*aG�%�\����� �:,�.� ��.�˓�č6b[_öK�'& `D����'�>1��������&n8RF������]W\b���{�T��0�H��s=b�t�^�*��/�N�@���G�Y���B�K#�Jʵ���L���5�rn�$&?HwxT�F���Lw!��\37ܖ�X��� %&�Qt���	[�7�봐k9L�#����pvyt!+^SE�X��i��4��e� ��;&g&�S��]��<rL˼ʪ�c�l�����]�R(��|>�o�sGu���p�8�H�?�FR��+�籕\�ykB��I�M�Z6��gP��ن��-� ��i�7Y��/�Z������ >���WD���O�=ԙ�^I\��w0���F��ce�����J9����_r�#����s
�CPH����Ͱxj�a�n��j1�:����<�V�]�ޤ|��A�,�4�c�rh�J�l�>�RS =;�Kq�(L��c�&�H���[�wF�����H]�k�r��Kb����nή�t�fq������7���W�.ӏ�>Q�Z{�3e����YВ3�E�:�D���<ϕ��¼��Wf�n�����+k
���0��D#I��D��(���l��=������8;j��7<6��B�wF����8� "@��.2�y�]���ч_n��� ��w���Ғ�b�5w@�қ^� �dQ��u�����#tc���J@�2�}��-��}���u�����O�5���'�����<��]̼��H�;�	��{d"�#�9)B[���4����ȱ�x�m��}��Z.�Z�)Q�i��m��#���jp�Nt`��������2^X���~�#82�R�WDAj(:�:����[V����b��U����4�'��m��َ������(8��0�� �+��z�q���~#Fr���S|������(P_#�vxjm�r	,��E�Ό:6n����l<#E���9w�b��/�|Mf=_p�f �U�L����La�~���ay�y]X��3e�j�������]�{�#���7�F�tk�@a���}K�*) �)|Xgr�鷻�/>ù�*�'p<'�ߧn`� 5�4₝5����bVFa�tĿ_/�����M�=�: �C�������� �AW;�~&����awNq^���2x�s2�O��?H$-M:e�z %�����"xz�ndy@�+����T�4��NeW�r���{[g�F���7GX1ۤG�7�Έܛ7	X<��hj�� 3R'�D���$���8ĳ(8�|7nk2�	��z���@/q�?(H�&%���aRj� ��� �j���oSTc�������s�_Í\2���qF� gqu�]��#��j�o�]|��H5֬�q��縅����t0Y4�9&����Ѱ�g�&J���f���X�4_���3j�ΎE��i����ku���ǟ��Mi��y↮<�Af�U��'�V���'5�K#˳/��|I̘N��]�!_�:%Ơ��=	���T�q��a՞̽���d�j�����S}߯���[�t����[S$�f���d`�ޅ��x�nռЄ���8�5�$Fg����i�_�W��v3��?�35�ԉ�z�C�N��H�HF������KQ�{0kHL���A֢0=�f��NŮ�J8<��;���Ra�v�]Av�/�BW-ܚLH���%"B�SS�Y�
���&��d-^(�z�9חfq7ѮhZ*8���i�[𶏓�@��hǺc1�����C�%^S��L=M��(�ԴZo)1����xDZf�4�v.��B��+�e�Dt D��h,	aS���NƲ�����]D�͟'��'�[3VJN��P�v�{���zS�W�
Me�܇Mɮ�,�2v��Ӳ�S�g�q���^���}�p���ɶ`��>�;�m-��8D�)����� y(vi�TO'2���X�!�!<� ��C`�0v ['uҜX�U�-ӿ��y_-&���!V���/�F��eN(�~���eEt�x��0I�(�&w6�9(~��x�w�{�����'���g/򮝝���)c�c�<N`y!��$��
Q\�t\�U��F���i�{]�s��HH&�<�Am�J�9��s��8F�R�����)������ S�h�v�C;pKTAڡ� ��w��`(?dB?ؿ�-���<m�����S��ZC���g:~��{�P9ﬦs�[��e饺�'j�|����"�c�G�[w�sO��yp���?Ý�� �Y>�jeQlQ�|��d'[�����`{�>����g(2@����P�̧N�R���g�r�Ik�f'���u�ޖc��	���ʸ⊾"��&uFhd�S_�g+ ?F=�	�x���n���F�{Tt{v;�0�v�}GP�]{� #���Cy�������^t�7�7�izG�)�ˈ��uG��@��_j�.A�>���A�s���@
�(`�r`ϊ)/n�WtњR�z��	�SՆ D�9�;H3袓�c%4
��/g�I��8j[��e2��Yǔ���]E�+��Ɯ9�ܙ.La�x�&aw��al�6�r���C����&���������*;$�Y�l"`�m�ǘ��n��P:���n�^��.�k�9nf�K>�Ne���Fw� ]k�"�V�2�g���A�&r2������z�4V��?����R�&SS�i�q�63�L䜓Z���}OX�$AE�M��v��a���1ߞ֣L��9�9�$���~Z��4'��,������C���fWu���؍�ևft��=|��f[�N���ǭ=U�^��:��7ʕ�#D6�W�@n"C����f���5ق�Z
�6�_=$�7'4Y����$�@��@�+D�$�pԷ���e�R�HVG������{C���tڂ,����ܒ�VC
�p��a�&:�U��4�O �E~��7�1)<��v�p����׊���O;�)S�Ì�%XtC܂���׀�U���\o�qm���T�N)��;)T�:� 4ou?=�;���+2�o���.�bi	����������8Q�7c�r���*�ٓ�E���|ӈG���V�����Y�G�2g�������f���[� ��z�H��?�2��׮%_]�OF�cBó@u�T7$8�,��(��#�Xg���&Y���R�� n�dz���=j�Ѐ~�S����K�����z�>"Kxג1�6"�q��s��"PVW*�7>�] �kaN��Z��d(��{ujH����F���m{�P\ਈH�qh�Γ��7�.`��~R>́��~�D�k�^T���c|q�#$X/�f����2�� u0��a��?�VB������bz�m0����E �T��GϥSM��Q���A��.��g;��g�R7�8�/�(��1VBF�Pt�EsZP4��'����__�
\�	���i\c�K;%�>���¡pe��p(�d��s=�N�e�6\���o�
�����rH�Α�������8�[r n����<R/��*����&tD����	��B=���W�9��.���P{y��������^���ц���U��ZSL�R�i��������,�w��N����w	zn�Q�9/�a2�(���$wB(g�i�K����>Pv�BJ��4�����ך�[��#o����^����4��j#�\��{�ep���>�¬e�H��~�&����ο܇�$'QV�x�YVB��.�*V]�������(G�,GP-!*r�9g~��R�r�?�� 9�IƉ�+jٷ�����L���0)�ݍ�X���AJ0Y]N$iX+�ܶ��+��e�[���^��f� f�>S��>?�m�f����)�j������In1By�k'�N��� �%�L��� ���>��6���y��~Ė@�����@�,p�"�"��=5�b���J�L#�b��;ʫ:�1�����ˊ�G@;�y8�uD5	���Wh����;��=�檈�+��
	ν�M2��m�b�=�P;���`2)�.D�'@2���M�ikftin�Ξ�s|
0����G��"���M�����֎4��K�����ٟnt���{X8��&��8l~�W��#܏Ӱ�� �����lݝx��I���<lZ/��t�Sb�']���`���� �j##O\w�ck�|ZC�u�I����%eQ��ɮ�z=��nI�\ٸױ(j��|�iܚ��F"���f���C��Yꆵ�h}�v�Ҟ�^����D�7l	��+vI �)�oh�q�������Q��"�7�~%؝UV�su(���U�ǂ?_�0����x��*-�U3W�*���%�&G�iV�w39V\�;d'i�����i���TD3�̷+�s��%�B}c����Jo��UG�?������Ł���������W�(	�6��G*����-�]ԉ���,̪��ixމ��tbN���/V?n������w�W�(�������h��O�������e(ө��ӿ�qͅlH�vӖ_f�����G�{��޸!������n����a
�2�!b0�d�(�f7<�2"�X�P>�����Tg3���S���֔�b�Jul0����e�!��+�(��%��d}��:-��Un�Q��4�����G�iKN����=�Em#�����[��wCc	�vNH��!o!�Mr��k��QJvrȡO����/P�!O���Tʕp��P>X�<��)�!|�/������K�l��u�V��ٕ�g�W������X;٪`���]wqd��&}HT�m��&I�2gq�Ƿ�f���Y+�W(~�x �+$�Ob��erN��g�3�pe6�y�����19;���o�r�^?�2mu�L��[�F�\2��Hn�� �t�6�R�i�K��E7�'�w%�Q�َ�А�Xkf���9Z����|�J�����B0�p�����,U�\d�-6�0�Q��C�j:��7yc!H�]Z*h����c	�$���/\��~����\�}�ֳ�t�����r�Zk�uxI����<�,��Uk �p��u���G����+Ew�ౣ�](+ߞI���jFD����^/湜�s61�&�A��(-k�8i9U����_��1���K`������=�9ʱ��?�ڴ=�uW&%��L5�D"Y��SS^(�>Z�C"꫎���;�{cף�)�Qb��Y�0n��>I���||ߋ����n���y|:ѡ���ǔf�h�+�����m������� ��o�y����4�O
��K��H�z'}�S����t��>�Ke�5�5v#q�Z	�)m��T�|!�x�0�m��0\�Kbr|i������لs����(c^�T�o��+n�爰q��^S�a��Hk����W.L<�PR���#�K?�d�"!����֮	�����K�� {K8�����Mʛ~���6�f�^A���ˣ�� ��?Q�W�)�d�<�'C���y���2܇s���=9�>V�}E��w����H����v�PS-��@ϝZ`S"�M]/[�w40��`��M���3`k�L�S�˷[&H����xzR�$u��X�:K�;��ѱ�P�@��5�⪩h���3i_i��bh
��s���lk�����@�1�����8y�W
|��2йBn]����G��N��$>70��X?	��w��� �N
��	�4����^q�ss����ݫ�SǿȌr������z����P�	��]��1�9��2k�����E讵�$�]���)d
3Τ� s���lA& �oՖ}�P��$1
�0�cp��؇��DG��ы���{�.%e�k';�&�-���,�k�DA�$0e���<�v����sp�2�
���O��m��v�H�,��R��}�Zk�y��ɔ��~�p!x�4�2=�\vr�.����J)dTDqu y�Ӻ|�9�]cı@^�/x�qkս�tݫkY�\���)��R����'c�rG�}�	�l&�Ό(�΀ӱ�h�Jě�t�y	G�aN�����T���v���딠U���	i�����P���m���Ƙ5v+d�O=�(1�{�vhɝ�b2������L8��i�	�lAh�M�.��ɽ�P�_㑩��]�{��{\�6!Ӣ�C355���9����a(q�uEL2�^Z�@d\������~�B�E\�[G[��XIG��&��S+Zɴ8�ߦ½�m�rY�/V �|"��6��pJt[j~��]==v�gҰ@eΥ���Ow�Hi�s�Mh�b�1���i��Q$|(3F|1�$WҀG�z���uV5��r*b�ލ[��8���mt98�_�f�=��P"��1��zE �0w�ma�\o�e�XjS�����iԟ�A�4*�����JR�{����M���\&�ߐQ;��H���C�!X�燡/2.�V�h%Og����nd2H��懒���n]w"{��Ⱦ}k� ?�Ȯd:�B��d��Y.�êT�5֋I[�,���X��{��E�"S�\+��QAtf�$���X)�؊���F�`.��T�Ǘ��(��f��o�~6�J��2 �����w#!Z�O�5ݠ	���#� �}�RDf>�L��5�e�	+6tR�_ךv����L˯v�P�!;*���o�l��:�$�����H�c��������^Z�.S�~0��>����r��!&�C�����#��U�/2֭5(to����f=&-�3�b���Y�.J�P��埡�N�W�U����8VBr�i��xgi�R9Xc��`�ca/iA�K4L�t�)Z+H������)�*4��zh ��'��;2	���q�>F�rmz�.�N�N��+�^�G���ŖT�of�|{s��2;���OV��m�G�N��5*rL��Oٞ�0�t�.
�L"y��}�U(F� ������s��X�p]L���`N@CW
�n�����H�'4%�蓰j�D]��Y���b��L�1!�p!�p���ֿ�%*���M�48hE����I��y@�'d���}tF�)����c�ī<��)�Y_��uC拓d�?>��A�,���c��ʏe�W�\�+����8m;��&���֌pl���9S���/��6�hQ��2J�e�}�W)@>i�#[��w�ǽANl|�u��`+2�
����ah}��S���yA��dHE|*�,�D��&#��T�^��`g�H��#�hi�R��I�ks�c�M��ڂ.�߼Vt�.�@��p����6�@Q����l�u��˥ �»��ed1��?%n;[>ZzS�����a��1�� ���9$��J�5hԐ�H���ӓTS�o]�Z3��g�m��R�4_�e��N���w)
w��ݲ1m0��pj�J���X���)l�!rv��j��v?D�����d�>j ��f�Yr�`��A�����;47�k 
[DZ�3�RV��h���P����ж�kFK��e���
U�����M�/��gsR-/��;H����?޽��d��l�<�"-ϊ`֬S�>`F�3�J:�!D��A�E�\� p� �)��y�sm�k��!�飶��ᓎ�>�
HhZI�v�Y�D��ͬ-y�d�O&�hͶ��ck;���C䋲!�ִ#[��4O�h��q�\����V¡��ݮ��Ll�dk+�o�7)ofM���U��d5�;�������gw�kz����4��W=̄8��; �*S�������eʣE
�	���P�kR,q��a�f���-�<Ѯ�L��O��ϛ,����z|F�֡\���V ��L]Z���R��Nخ�e1��×P���1��I�Nv�E��4-����M_Q�Ǒ�wb��0��T�סt�׋M`�an6��ׁ�nba���0#+=�|��|��ڐn�Li"�,�/ �V�yxްp�{,�,Jح0��|�`Q	�摱&�ּ8'��X��3é�,���O"��&��]�?q[VYq�k�� dڝ$L2�5-���$ӓ̀Ќ>>�����p&U@������h5?)��q���҈�<�����2�	e�ۀw�VW����J� ���i�z�CK�*ӞgF@���L�@�ι����oF����b׃\�ȱ��%@��R@�:fY[/���}��~m��Z�p��e�a��tLa< po]����7t��I�����lZo���K@o��@�!�Tl@kEނij�)d��?�3Uy����W�}E����)�@@X{/h��@+5],I�d_^��_~����2uj�k^�i�u���Uj|�h[2�6j>:Ho-���4y��<��[���LE�X�]�ЧӢ�Ԍ]2�XFD�3����V�~�mm7�YKG)���������<�SۙY^/2�nU��x�Ccl�r��m�(zn1 �^.����_�|�D�uhd�T7�x�n�ulVg����8Ɍ��2��̸�?G�Wz�F�pL����ZN��~�4/'K��K���\7<̯h�Or�p3(~��G�a�Ǔ����燮��N	���9(�U�r�	���ܝ�"�Ɔ|��?�NCat��f�R2�9T�d����+���)�mQ�Ry�E�a�1l3�sht_�&S?�g��l��jc�$(���)�N�G��뾮��9�����'0���h�����mתS ��6�!7���6�6g�w��J�1E�5%� ����U(��!$̎�6��Y�d'i��-5γ �ŉ�!����{
����D����냋�����w�����C�7�_���@S?u|�� �V8���@�0*��/�g�A�s�0�7�� �x,�
�̯^�ۡ8�si{����=��S6
��u���P8�h��5��ϝV� �hAڵ�A���P���%� "�.�C�`���1(gIl?	���	���"���e�(��]��X�K�a0�*�aA#x�Z�^��N�0u�q��My~���8�<���ov��Ol�G\��Y�| �~p%D׵)�dW��D���XG�Gp������7hR�������Ñ�b%�K�[�*֟�;n*�B�q�}8hx,�^�� ̆?�@�2˵͘��Af�~�������%�tY}"o�Km hkrbb��禲��$x��T������	������2(ң���I|t�.����.͵�gV��j;�cK�'^*��(MQ��s7�7�`��Ὰ~k�<���Q��9�\S���3�eG��"x势�	�ܪ�^`�K�@K�D	�����@�P��"�$U;�n���w�&M�!T�hf��NW�¡�'���	3��yK%QD�5������!ـ�/�t��s@%��6�ϛ�#e 3��K�'�2��U���D{�-^�'�n{fkv"ԛ�ݝ;�Y�	�A��`���p�1	� �[#������z0�Y��w�(`-樰�H"��\��,|�7qo:l"&��Й��fR.�����Ju�b�6b�s���{�UD( ��Ov>d�|^�v?� �zr�eJl7v7~(� 2nw֧+y�>�d��Yj����sBRs�{J�O66Su�Դ��6z%��lxm3� ����ܷ��a��l�a��U�@�}{&Ƈ!�EQ��-����rz��n����>+����(Bb�b�j}]��
'8i�����H��d�5ƲN-�����)l ��3�X�� 0�~X	(�apNzG9~����Wvn���b�ڝ�^RB|�\z�h�n�~�rJ~)c�����]���gm��KURE�����`�2�)�`�������^D��U^h>�LA]�ߙ��BN@�u�۹�h�%�?�9�$u3 �v"b�R�^�p2���)P�؋^VΫy�Ȋ�4��?k@���o�RYĀ��~�Kύ���3���n�yfۡyH���&���j)9¬I���{w#"�:(��%� g�b?�:���U�S�<�$�<?9r����eܰn쮨��]B�j�K+�d �d����S=5��2DnB���7x	��~|�͐�ڹ�)�|����0�X{�+�A)a���W��|�U2��Pv��rQ�Y�=YN�49{w��%���z#5�l�j}�S^��?T;u��M~��s��1Ŗ4�M�#�)�}�{x�Gu��9c��Q;)�f���{'��e���J���wIp��~��u=?�K���Kn�K���?1IB�m���R��gz��7��D��1�S�����J�ߨF4��C'��ۡ�%D� ��<�a���)���am�[aA:5w��J���^��:#�V~mW��p���ڲ�.p6���xZ���T�B�5�|/����k���Y�Eb�jAW0�2?��z�'Z�i��IRB�VSB�%�$C5&�2�i��df�I4�}��^����՛CXd��F���@��G7�����ŗ�|���3��%�v��%0A�a�
 �W�g�m��g3R3�z��zl��s����ĉߖ�<})$�7ԍ�e����VVH�=����v�1f�U�R�m���S�=!K�c�rxR�*dЌ+�Aq҄?�6���7�L��v�3��(u��[�'�gW�뛏g�3q�o*q�R~�~,b.��5R{I�W�A�Y�H�q�1�'H.�E3��qL��������`>Y����|g�Ն��{r���$����j�&?�i���'�
E�y5U��{��1�A��j�~*xW�[mq�a$#��Dč �s������a���� %g'G��\8�C%/
� T9�;5xK �Ř�ބ����r{��w�8s�[�^��%+��J�l~�t��8H�2=yd=�~<�&�����B\���o����W)��zcp����Qn�#jFl1�@8�����.,�I�/1g���F���D4n���M�$��~0L�A�ɩ�Knzx�Xx�ʁ�X7�O�<ڹ��K�m�!OL(�����Lo"M�}�g����� u���2���$��tQ�.��Q�����FG�낪�$Hѫr�$A��i�CIb���\����^�L"�@H\ȱkU�@�������U
��R�x�R?eރ*�8ra-��#�3�Ƥ['$�C�후�n1���a�1�?��u�w��}���>/���q�E��~�Y7��U�;���߭�j#�vvem�jaQj@��|���_tiB�kEɬ��������/�7ߛ(���M��s�z�<�"����Vܫ|l����X�Jk0����s��1Y{~���a����}���j9��[S*����z��զ��WU�S�,�3?�CG�ߖ�!|�,�ć�z���yk�N��y���z���y޳}&|�Z8Sg����D���%�2�Kqa/;�<i�ج�.���*Sh�Hy�y|�P���� �������IZHL�'Y�}��X0�:j��D�,}���I1�������WT��7|+B	�#{y0VËK��(��w�x��|^��͍$�IIsQ
��`FI�>�]o38��&�h^~�i��m����������SQ��y*#
�&y��#6�J�M�!�1v���B[�/s�%
�9�nqP���6@k�����_��96�Q���Czai┆m38f�hԻ_�{Jѭ|����a�V������r' N��U]Dz�I	((7ыd���!3���Q�8-�O��V6�������JU��vUL8���[���T�`x�ڀZ��
�}�'�h�5R8���:���apOIO�^ u��H@�ޗ;�̲[����/9&�L�lEs�8�S�����}%_���BLa��p����S?B'�A)&�j5zރ#�_���H��a�~xF�xHUɣ%(ۧ��l"j ��r�(!^i������-��SϺ+u���tyA͉�Dlr�8�Q��]u���=e'�X3�,
��A�F��׼���|.bLT��)UN�dPigó�N�D$�2"��̠:�Y��a��v�r�{݀g�?1�"2;�������������<JW��⫖V����%o��@�9���4
���V�����;^�76�)�Y�3{g��5p�"�9G�-��?Zf�js5?����U	~�i*Բ�Qo	n��������n�^Z���������	&���C��~�i�j���Dcd_�0�*��b(�T��16��81�&�����5:��p�t?	�Ah��#�ԣ� j��{�,�d��19��5�]��ln��\8!��oY�4�k��*;|�Z�ugϵ-!@�G���XmaB2c�N	���m#�
��'ݳ�]�w�<�є�+ND�-�+9w]ZnchǥwG����H�A��uݗa�&����%������~���#��ur�8.��2Ւ'�'tT\5�W�"&�Y ă��Z	�*�c;x�\��T�5�#2�ӭ�\�8Jx��p@�����ڍزJ�p�eR�˧�R����U�,�g<}[3�M�h[0���ʝ�KA��#}���aT�hS,�DR)&.��kd��Of�
K���b�+X)^��f.<�h �Oi&h���u��c)�_'&Om/o��P�Ƨ�������17��&�߰e,�W��e^�O�a=����ĥ������<�� ����x�\������h�b�Y�E��O�p�^�i�P��^���0۰J3?"�W��S~	)�<GQ�H7lp��m4�j�Q��Q	��Zu��%U��I*��á������-��R~�4E4�z�I y�1\
U��8I�t����w�'T#����|�.&���-�1��Q���{oNS��|�ޛ�eA~��q��<���毬��Z)*��Ӳ|�� �(t���s�w���Oa�:�;V��/$ZnN�Wm���i]����T8 '㋆���ء9��.�R��$'���٧�o_;�a�m���lǷ�~��XfM��v9�;N\;�'��'��z���[�法Jl�.;�L�yD8^�P(�|G�:?� �G���.�����~�
\��)G�n����f�td��\ଔ&�O�� ���O��w�)fdnQ���j)Q���GHZ�*.e��gw8J1p���\�n��vcFN�B���}f��6����Z�7a�yK����
�̸[�B�(v	�3B�ȗo�ĩؼt�*�4,"�@O�=��a����6�,`��V�T�R���&B^�1�afq-�ފ6�8I��]�Ì�,�Y���Y�
y��JuY��^p�C���y4o�pM7h�!�v��.'�gJ�Ny��|s�K��L~k�W��ߓ�[5�uD�)�Ҿ��U"�$z�w%??̶?���	�ZZ�)T���$۬܈[=��p�	7ah��5:p��wT�P�}q�Fs�*C@���d�U��#�u��<c��p�U���b����c�����B�2E!6����quoG�:)�.�����Z�e$�]#9$g�-�_A�Q��2:n~k��O��|'㺢��>/w�Od�q
��Ƅ+�lߒb>��@��8���x��co�?Q2�L�����!Yª��wu����Y��1}�I>��zT]��P�Y��Glr����?&��H�Ց���`TڤԘ���/^9��C�A?M:�Ü@�X'��{s�6�P���j��
͈�4� >i����QZ�K�����E��|2����0Ԉ�}�Ųk��aB9y#�_�N!7'ʝ��o8k�+����-�	��h�iR�$�!
�pv[�ŏ��W	@��2x\�x��+��_`Գ�4�H�5�T	D *�82*3�djR8��c]�)8V{�D���M��qL�Gj5dF�;dcu�>�H���A�
i6{i��A�y,�`�O򃘏T�����"Um�ss�[ް~i>W���Vd�4�@�R���r�u�c��CS������[܃��z�E�F���YM��l��^w�~95z-�*��K=��!m�v#pl��u���UP�r����EM��\�w �`ﬃ!��x���{EHjK�i�Wg �E�@9��r�,����C��dq�4۝uBw�l� g˭�&N�Xp�$�؍�EP��Q)��y����>�8LҔY	�S0����B^�Q%h֘YO.���*X�3��6�h�F|�� �Y��MfH�2�����'ʌס!��/��a��w�"�a�n�E�MAɭ��{Z�5�����H��S�4Ǻ7���K��/�d�	̋�ۙ�w��F΀Yǳ+~���,����FLzϰ*��N�\��O���)�:S�9xoBz���y�VD�cp`4k{�p K`�g��5Z��.��D��Y7�D=�oz*�~yTBX�>�I9�����7�O��+�a�EB��\Q��'��� �wn�"*��A*�>� �S����OxT����N�#�\�c$���f,He3��MF>^���PY���2�lI�������e����-�\H�l���$yMꄋ!�ƙ 2n��no� �\���n�������0�D4�Ѝ@�ǃF��P���o�C�C..������])��1��)�Ш������c8w�	ws]rA��t=�>~[E�;��j�� H����g]K]ЖA无�,h_
p��b�YWwH���帓�\�z�&�~�6��O�\�Q,��!��<�ı��:{1Qw �|��G[>�����.�e�.��)5{���!u��8R�	�9��y��[u�-R
���)Fztl`O5\z8U
��mN}d��23+uɠ0zn�'�U=\�)�rL�_WG��\()�Ь���[$QĻ&�!^�,��{2Q[����+��Aj�����Ȩ2��KvQ��nO�v�m��tխ��l��L�\���킅Q�(��o�F�иf!��N��A��e�W���.z�:qӑ��uk��U��g+�~u��4�<��Wc�C��z>�F�(��ݒs��.C_ �Zh����s�s
6�ń��)��b�x�FO���X�e���a������A�� ��X�4L�LJ�UCa�e}<v�.r�b�9>PL=�}Q֣��azc5��{mN&��¤�Ym������x=�R��$�t���:�g�i��)��T�q�b"�{Xx�r�׵C� �r���_>G�d�X4��$��f��f�S[���W��O����v����ß��z������C�P��:�.`��b6�,�-���h�34��H{Y"�a�HnE��(�*gDݛ���av�FzI������+�w��7��;ɨ�� )4�B�M۠�Q�:mU�Z������<S-@#4��u�C�k0�����u�쿛h������ѩ�,���w��e��q��玙&oY�w�O*�m�U��Y�4$�	qD�H�Xe%��K���~�&Z�����	;E����?R䁽���٠&6����E�+V�y{�:won�0h�q�j�������>!�@g-��W��M�������Ա������M5?=�L�7E�/�a�`I5����zѴqsy�w�5�+�{y�>��m�0�lR&-�d]@I��u���;�/S~'���V�5�A��q.9Wִ|���t�`���!ۣE�I���(��ȴ��;�E�,|��pM����m�I�F��r
�b��*d󉀣�*�C���݈N�!;��E�~l6�R�o�,:X��SCB�Yw�ƺ���Y��Y=v����۝�m���	G��%��C �����$��(v��a+�n���`��ʛp�������J��飲[�qf�ἱ��N��5��V�D��v�C�ӆ�7\���s�މ͂�azE��Hb�>��07PV�[�������T��X���(�8�7�%;�e+:�N�7�����> �����E-M=V���sr!�Gǖ��)k�{Yjs>�BX4I��MqJ��1̣�Ů/S�r��
�X���q�-�տ��F�b��%�,������5��E�� ܻ3l�U��R8A�{ScP�F���3������T���b?�
O�K��r�BN\s۴-2��f�;��7H�S8����Z6�n6
���:fo����tC��r���@��S&	��Y��bՙ;�T̃�� �,�D����xԈR{b��J:�A{�&�'"�0#g��\���ͮ)b�̆�����ϔ:������؛񭾱:>�9�̦������������+���x�z��i���*n۟甡���FF�����az~�U�}��?X��i�vM���{<����*Q'z�i�\-vY�6�&���Iry��x+�	��_`"#�..K/}��ĕ8Z������[&I�7P��R۠A��Muf\T�Hx"3s��x�5�@������E)�����T
���J�N�U�d-cmuL�4�jG5G[� w~Ι��tyW�I@;��
�h�3�IT"�7?������ToĈ�W1�d�<S����e����I��i���Kt:��FF�~c/��+A�y�C�;_9� ����b���y�y{y�r�U�]@)�T������|(kBú����i�r?RM�9|�Z��j��;���i��Z�����C��5���z�UvB�{��zꬩI�Ao��kXľ�9!~.z�\봈mSf~��dps��K��ޖ�Xf�~V�ȸA�"�75Y���!�F��㆞t'��y���s+�m�kB�<��Is^��m#�l��H�郉�x�	�u����W�^b��=��Ws�"e}��T�n|�fo���E�	z݀���D���������}���_V�&���R�l����PU�:6|�v��9Vz���ss�`[Q^�j�ޣ��+�?zB���j���첉����?CL��腈�~90��Z-J�^�9����h�8Sfo�=�TS�nx�v�����1#۴7#�l�T[:
�i�x��
�^��!��gEW��#�K(-�tj�fF�e��uS���΄2he�Լ�T���v��?O�9�@�G{"\�*�s*�j��x�Y�Yd�A�3�wH�ҵޔhj�_He�3�� �p|�˕?X:~�WP���c�?����(�ڲ�Ay�P�
�E1)��!3�\w�$���K&�	Q_����7�����Ht�@&V��S}�u间 ��Q�)Xs�y	�T���;�������u��v���5�p�L��`_���!��=� qCDs1O��b:]��׍�f��?hN.�W�Z͚I�3��O��N��h�k3x���Ѱ�a��,E(����ݍ���j�L���0~b�.�����dD�*��H��n��K~0�����.M�&��^���,��A9\݌ [��`���\��u�f�q�M��-���*�����&�<��ɲ�x��}��!\$�<|=1��זD2Ԏ����������Ū"���x��^Y���ԭe1"'��x/R,W�7!�ն����ݔ���ăz�`9lĹ�9"����������ipI��@: ��w�C�^��;�Gh�DQxT`��Ծ��X�4���n*!/�:�d���#��_�0߬�!�T�6�I�;`経��_P������ÆX����җ�z����y���TKR5�S�����6��(NԱ�u��!��c�x0b�MG�j�4�3� 9�>���J�<ӖL��)�]+����<Ƽ���Z��l�z�{�*�W���pv
�)3h�iݭ��i/b˷yrٵ�t��v�=/l�\S-�0�vV);j��7�(4o>Az�E��I�wY��D5p\����o���O�"�˛�=>�$��:,'T
^v���8���.���U��gFJA��b�8��]-aHrٷ�v��/�ȍ�b��H���b3�p<�]�f�H{XӺF�a��"T�Ii�%L.Q����^���\�o�΂�a��4��R݌��rP$��H�����j������ �M�G��� ����r���_�Q�2�j�O}��)��	�n:����i�ګ^ `>� T�����{��k�Oȴ�ȫ����?-�t ����w�fC��8��3vfH��ڰ��hX1����k�^�\˗�Ň�h\\�M*�E �dK�e�O���k�
�=������S��b�5,_ ���2/�Ⅻne��}���b�y��<n���SO{W1�M[ذS�r��)-S�L���wO8
6�-�ɱ�
JN������t,ڦ��I�����mZ'��E47��� ���Kj���FB����lD��8�J��ʢB[�bv��9^�vq�wdP��޾v�W@���y�6򮡢�U�]����e�&nX����ޔ����##54���?D�ư�@k̞H�&�39�=m�t���D=�?B^���%��v�Q z%�%b��/%������1��\��C�z�̊�*uu�G�_�rzu"�������'N%�J����";�9���s)^ND5���d��%1�x%����N�V=��P?;���*������A��$ݩ�ݱc��U�s^*u��ހR #�h=ƏZDh+Q��rF!��)�L��E-L @�>29��g�}E�Uf���1��/��.�GtF'E��������ni��=-�W��b��,��	n����<Ď��gC��̓^P���	�8hlG�>"&����dHզ��"��8��6gQ^֋1Z!k_����~\[��R���c84(�G�$���&ElV�v{5CU��#G�\}�����DP�YI�x��ԣ��aV.��lE�j\td�(5��T	E���]V� L���(��i'�'j��@��=ɛg��'M&ת��b��˂�/O6Y�L���a�]F�1-��n�,$�IF�HQ�B�/�����#�\�/��:O_:3M�Đ���pP��4$�O��hՏ���|�m@?WX�A	 ުI�Np�-�\qD��M�?�{�=�����d�3p�Đb�h��~fǯ�A�����.�t��ʧ(�^�=��l��@'�/Z������A�8r)˂����1�l��/�|�\ ��NX9��ɺ���\�y|�	��S6��A�<�	������e�\�rm"^�!Kk��!�}�!�|fՐ����&��M��&����Ͻ,�#-�����Q�:.��A�
�W���۟*ja�6^r�L��6��/�꿰7h�-����Mҹ'9���w���T
����:!<�@�ӵ)B\`�SK��Ģ�c�R+j�ך�;�R�����#�B�(���K�Z��*9jl���S�)�������?_�|�n��"si��\�:�<�yO]L�g��$2��j���̓��sHb.	�X�(�'@��?3Hv�������*k�H�y��裞�r �W-�$��~��4�f6UE�I'Gj��đg�N|�i֤1��B7^��f#�� �0/^Kp�Y^�mNWx���U���v���SI���B��X���t�m'����C���$P1	+�G-��l[QvJ.{3�dw�+IƆ�]P���&�,�e0�$��T!
G[enUb���7�z�#S�ю9,��b�]<�7�T�ByX���c�׻��(��H�>G����yK�G���_b��I8��я<F��ä��;��K���� ! #����5�wl�
�y!��f鶠^n=8#i۰BG, {˟B�B�ޤ-�X�k2}���C���s$�-=R�e�i���6H�N�ܱ'���d����(u	A9����"@O� �b������iW57��G�C�4	Q��������O�S#���ʆ�c�p���+`�w�`� �0��(I�,?��Lx�.";�+_*�;�&O\�HZ��?@����&�]�(��]�y&�� ��:A%�>%����k.m�;�����23��R2I3���s��$#�)�د��+����xO��,*��P[��V�Ӈ V��% ��*9$���@M33�M���fߝ!���5���6�_���],�p~
H�(-���2�Bq1�3��~�K��Gx�D^���v3�C	��OH^�c��CI��#��8 .��/-y��"�2����r��2a��o�BM*HKf����T�g&���Q�.t���h"�jfL�@S1��s>-����gg�
�,/��с ��h�zj��u�ޗ��ƥD;�Y���;��� ;��G�{)\+}@���Z������"W��>�KݑrB�x����(h
�PP���'Rse?D�V�6�fW�#5+v��X�V"��d��6��Y��
��G��.�^���w�Ź�P��?���������q����/�������-��D2��hɇ�a�wV��P�}{:DI�{�M�"�]��:��LS����9}"�v���|�z8N�Q�e�~P߈y�IEM9:���0=��]��X�ʒp^���b��@�*w[�(��NTR;��W[�\̜�$��-��lݠƐJu���'�� S@",Cz'�S6�k<�m9^�"7���9��賰[���`R"�Т�\?1�����J��+�5������>M�,.�q�* V���p�w�g���N�*�M�wN�BÛ�����`M|�pkT��U�VGLBE��B��f�
s���hM[f�qL��	B�R4E�����J�d(����A�w��ʬ|��N��/0��/X*ϣ��XY�����{���Y�}������t�D�y)����|)(ԋ7]�|c3M�_]9%6vٍ�hK5�@���kddyhR���!�-SN���Ǖ0��[�:$����a�G�N��mc�6��8��|�5Z�욳�y-:���`�&.�t��	m�1����>K��y������t2*��9��P�az��.��z�=�Až��c8����+\ת]N�ݮ�5�g/��<|�-U��-z�;���]u-џqm��J�U���r�!V���x�i�S�̝2�	�F���\�h�?���]{mB#��|�~�q�GP��ߝ8v�5LxxV��I������7TG5"���C�M��/��ț�:2��*���|����5D��4 ��]�w�B1c��W�͛��{V����އ��+�i!A��ȁ�7�C��`
4sʺ���VE�j�vw�٧�:��o��?�7	P�����U0��1�:j��"�H Z��^ٲ[o3w�Ka <�%3��f��$��"�Rh�k�fDV�^ ;�jW�&'a��&���K7���-԰;@_aU��E`<=ҬY�p��F�ʸc$���5��rX�����*��6����GҐ�������yqT$Yc ;���Bc���׽ljW�h��{T)|B�� ��]YǓ#D�>��"8ڿ����I�p�FU��еn�N���n-#\O{RT%�kN���hH���ק�{�[��ٓf�{�_!>#�a�Ľ��Q�M��qAbu���?x�	��z����Jv|�(3����>z���P����&��c�3.>Km�黱�NB%w��sT��8���~amf! 6K�O�؝�����,���!o��c^>�#�l��B� 4�0����v�"�2��z���|�I�(�8%ƶ�@2!���)P8oC[��{�1'����o�J2i���{'�䄶))(��$�|�8y��!�ӾM��į<����������xF[a�+�M�O`
G�R��w��3o"m/;K4f�n��nPG�l��4R�u���d� �I�3x�z3�Q��'�)Su�m�/z�9�f�~��F�p.L�=!�Ex(��g����|���/�)�bX�=�0�u���D+����y.A]�����y�qgh����0���# a�D�4d8kS�o���J��@<,��.�ȮVI�d�x\�������O��]>i��!Y��o(7-�iP�eׯ°����d�ib��[�x�k��(I@�*2�TF�%�y�`b�+�fS�k��,Ih��՝k��
 3ų=-/v��xxHy�x7J)廀y>aHO��m�2z�������`��a��o�8q�@����J:����J�����VF��)ʹ�S��g^��n�r��5MVO�,.O���3Z�3i�_S����n��M�P������/p���j3����r�h>���B���p۽<����{�_�����6D�xlMwi�b�VP�S4vL����<ѝff�Ӵؕ�A�_7ѧw�5,#�Q��tf�0t�+(0�����ث�v��kX��j�r�'e�Z(����2쁣�����?vI��iӿ>��&Z���]���r�r������>=��C�b]p�â�O����H�-�|��O��f^N��s�6�~�<~�c�k��hml
���~���)�B�5�[�+c�z��`���Eض$!G�o4�}��;5�l�'�ⅯL�B7�m�yZQf�E�
�^�<(w�$�H6��*��Ƿ[� ��^�JnO���9�nzb��G�
�eG�rOd�g��}�:�l)�&��W:���zEKx���-*d�Z�KO�ߘ��	''���+3��E��lM�+���-�	��[�c��S�{���+;g�o^0O�UD��?"A�I�k�_έP�F�ԛ�;w"A`��ؽ�-�%i7�z�(��'l�I~@Jk>��m�.M�5Hi]�'��/�N{{����G���x�akDb8�%��"��Y�U�+������ǳ�Y��#���E�y�I�[�7\M�'y)�:w��F����A7�E�u5d+:��?h]A��]s��HAM1�8)�`A��pn���P.�I2zcy;����_Z�d����*]��vX�������v���ܛD?�g�7N�g���aWR0-%�Ç�hK��~7$��O��X�~`�uo��2g�FA�(]�x��nq�M�ϯ]X�]�A�����DW�h�TkR�ü�7A��g�T��j�1�Ǆo9�������U�ښ�#!��v�qz�۹��S�I�Ջ�Mq%j�c���^ys5�F����\��\�S�){�d,���*���0cd��Z�����X%������n.�#}`���xZ�g�w�j�f�v�"S�3���oC������	~s��ą����U��^a7���7��\�]�-��MV��H�ь��m6�|�2�@^��|9�.�>��%�?M��Ơ�)�RW���\�U(
�)
:�WK��j�������p�=P�u�[�E���x,E2d�Xqi�Up�f��{O���u+덬�`j�y���kz)1�q�JPu$�"r .��)�.��&4�K��) �L�d5������W���]��6W��e0�����L����6IMq��6 b��^q_.<�Z�q%��Z5���]��~���K~_q���~Y�^�I�C8�u�3�� rL]`,�R�o��Y�� G�p [��P��ju��;�t>5Nb|��W$�i���q�^(VQ{N����؂���Tj�{fE^��Y@��<A�V�*���A��>f�>b�QE^y��xJO��8S�4��q��K��[�4���c��"�y!]m���c�e�S&���l%UO�ԋy+ �oz@��Y�1�����yL5�-|2���;�,[���	��>��˙�,��9�[T�l��^߀4��(I�L݂;��\�?�����7!���5x��Uc�rp�f
������`�/��1�Q왁:�vRP+����(����beJ���bS-�_��42��y�\_���k�2����&*����J��g��S����z�}I;V1�cw\+��d �R1���h���?�yX�r�!d��TA��u�Ǥ��b�SZx�����k�� �+E>�!�;�eѫ��12/�Q�{�E��e���3	�)r���3���n/����b/�O���BE����$Lx���2���3���Bv�P�r�\Ll�R+�kqۇ��*%@̑���[E�.�꫻�:�,�=ls��~w����6��.��[ sx+��5=7�?Or|Z��c���$X:�E!�lJ:),��:);F�5�����|��	�6jP4�D�����àl"��4����� ���LӅ���f�H%�D�85]C�����)�ggh��4qs7ܩs�o��b*Sn�zm���,m����Uz�D:v,QtIO�4���pGþ��{�ST|�)|4
���[lg�:$�Cn�+g��&� �n�ɷc ����D��Z����Gģ��lW?��wJIl��N��l�pU&<Sy4P	��A�b�`I����w���C��_\B��k�����"ʲ�7u��r݈t ��S�s�*� ��� �:��	�K6`����U��7|�ț��k;Plaȃ-h�;X��N�����a��[�D�E�$�����k��,]����u�"�l-�5��v}fh�(J-�g�����S� ��ӗ7CM�?.��$�Cf���L���V! ���U��pBW��$Oا�t���	̈��$�(0񤿯tKs�nv��%����6Oa0*�_{6q�H��au7v�%�؊[�С%��G���D�y��<E�`���0�w&�"��o�q42�P{�~vWѓIu�be�	���Ԃ���6J?:�#}����L\�&�:~��E����=/A��7TVe]W������Alo|P�7��ɩ�J)
+�O�3L12Jr��4s��0a�!�����Jr���a�Z�.�U� n�T�^%Y6�RYAr��/h�.SqZH6K�}$��M�J~ר�>�N��h�\y��	�0���/�Q?����q��&�o�����v����Įڍ(�����"c��Zb�y�Q?X�A��:�]]<�'5J���it_|pxO�OI�*P�z�(w��a��PB4*Z��(�L�/�C�s%��p��"^�B&qc���bל�bmZ����p}iB\: -n8����m6��A��BF���\e���nc2ԕ�����I|X~[y}+$^I����[�۱]�q����@ 6��,_�faWD`�t��S�X�h��V�ƾ�! �;�J���y�yzv~~�1����L����C�)�h�zn˚���ͼ��TZ*���7��B[�;�/z&��U0MK
�N�Ivx�`Q��\ԇ�6ͯ��~��e}R���$>=t0�E�pTb��#@���9���s����M.�_� �	}3iN�{�*؁h�l��HS���VEs�_^qF3>�0�^�R��yV�|1�yG��Wt�!��ؿ��n66҄?yz�V'R4P@�y� �>���}��C�8��n����h��]~�#�q?2�B��ث2���,�����+~�-
'i~�M	�����OJ9,����뉳�x;�Rx}�+j�C!��xB�G9Y�	NPn�b��jwܢ[$L�	o$��� �ٳ��Si�]�پ��U�7�_<_���/�O���� @8L՜~��3h���f槛�������f[<�h~T�|0��W��#��	��r5g�kWی��ŎΟ$�X�B�"���C���&d���f���|V�\5'1�J��Gv�f�{��?���[��A&��$iYs=���㠓�N
V�G����W�D�V[��Ð(��*�R�w-g^l�w&���\�-[Lxs��EF�@���o-fB^����
Hm�C�L��~�)����ގĭ袊`������w���;4�	7�ט��	Wc�'�T]mGGq	��}\�M���lz0d;W	�JEt>�/V
���Ҁg�{ր������ص����m�R�^��*Ĝ.������6�QZ%��-��(A�\t�/"��zp ?%o��8�p5�WU�#�'��|����kr���ZH��A�U���%���v���JYǫ�|�3Fڈ],x�w�;�\�=��]�-�HRL�8���a��P�x����n2n���x9Y�
�	 b`��l��R�x�o���kR�6�� ���S���=m1)��:��
�9�p�Bk�Чt�{{�gn��w��G���X_���{�kդ~t������r+��Gw�� I:K$��vㅇ9$�r�����x�O�E�	���=�L��z&�{���nr��������-xAdE��7�OqTd�:D� �9D�1�BrT���P�����������N�4�G潆�fݱmQ������H�!
�4�b�!_�%Ga�o�ؿ<��S]�sȶH�{_�D������@���vgj�K�ϴG©	��&\]Ew�����Z�1�k]�z�,�`���ܱS��A�y�(?�o��������A��cL�N�8�jユ �u'������C&�cj��|n7'��]!>�*�v�'�:���ـ�yѝ��$�[�qf[���O�;�\��@@���歔|���+2��L�T8t<�< ���8N(�r� j<fA$�DH����h��$���)���'��pHTG&�T9(�����L_�����gu�+�&��U��q�1�oZ���h��c��,�:�(�w���Z%Y��@zN��)�
{q�f�r�GY�`k^k�:�܎����G�d8�(�M�r����=�2җWᡋso7�i	#1죽R*�W*4Z��S�x�be��Ĵ�!�k����ʜ��,/IP�]�#�;E�٧O  wMXѹ=7,�v�Ì��P)~�οP��~���b��}�kA�q�R�Y`��r�K��'6��f��N<v��;�fgT**`˿�j��aݮ��!��Hp`j�L�s�> �I�cR�o�o�FѮџ���kј���ڢ/�ۖ�j;�~���S�b��C���Q+h��oS�`w]�*�,���G��<�O�@U?ӹ{g��YJ��tM�}�(��� �0��P5
�E�Vb��=TD�ۖ�ȣ�R��/�� ��n�&^�œ�S1(=s���~~�of��tæۤ�r�{%���I���_��,.�\PHnP:�$�:�E�OO��(�7ӂ���µ���9��C?�s����5�{�����[]��W��WD�ܷh��9 ~1������&h!;2*79��.�{nje}`L��R���/����9��ߤ_ͯF�^Q�IvXx�T3��0jG��i?��[�3�E��-�n�3k�ve��D�W岬s7m�&(�U«�Ж�l��m�RQi�St�ٙ/�xs���QQH(@ۃcS�Fj��c�&K��y�7��/7~E�,��G��?�0G�2T�x+%�<��n���';�����bT%��aKv���[<�s��K�k(o��� �ܲ��X��UEj��= 8B�FЮ�8=�ˊ3�]��;�#�T����5����Tox9�]�Kp�U��������B�GA���Ȩ����9�Bbk�/ P�=�H�¸�S�ZE�g�hh��z7uI=�<&�wp��]�O�Z���i��fx�o�	���AR��pæ����x��̍i�E�N%�*�E��(!\͐qN�G:�>R�m�P���$x���K#u��定R�5g�<l�b�_���Q1��2���O��W�葏�>R���v��E���W\��5e�0�t��E�] ��E�������cpm�5��C�����.
�4�c���"%ǅ-6���H;V��1	O�57��IS����.�ADzl�u�t��ܱx ǩg%K������k��j,��YX�}��ㄹq�����,�����9�f��iz��dG\�V�z#큄F�!&���7?�m���u�*:��d�ٙ��f��K:}���Љ��R�.��{UL�	ʪ��A��X}��J���.F_T�&2���sR��E}� K��(ݽ��m3�
�m!�Z�7b��i��F�N|-�?B�Ml����Ĩ�÷�T�V�|�E����`���T$����_�#��=�F����Q�a�d���^nz&�!�d ��1��"���^�i	M�+։�����\�T�_ʧ�6"WR��Qicsz/�̓>W������[o}��g�Z��[a7AU2���@A=?9M\�=@���Z9f��������4�H���I�|�
Jw��#�J-4�V(� ��1������!��YH6+N^M�o��>6]	Tٕa:-�k��Q𼇆܁z>���?������#U�\��9L|m�舗�W��v����؟7g3!�G�e��Ţ&��"��/JI��W*B�f�/!�B}j�G�r��Eu��9Z��4�6�~�rZ}�i_�S��:�
�%�Ơ��wP`y��..29�l
qZ5	.:�MRƤ$�*2��I�×�{x!�3�f���T�n5����4�e���ꂉ��~J���r����1o3����頽��ݦ�:�SA��
�����?������L	:�XCKP���V{J���U"�+ l���f"ڹ,(�_�e���G��	
����OJ� ��d��3A��-f�4����e���Ӥ�.ޞ?{5�FV�[?���4�ׄ�>l������b9�Ж�&�B]�jn]�9������1J��BM���Z�b=�Om��mC�b�<*W�.��>�R���Q(����S[����_��v���CL.��x0�Km6Ɖeu�ߚ�i�F�S���nG���{���ȓ�<�N���]�s�����2?��1�,-����ʘNő9�Ť��W�/= K!co���e�N�������Bn�@VW�[H8��#�q�v�*�X��7V ��.��P���T���+Z}X�/<�ͫ�|{=���W���o���F�p��t�	Q^3V
"v��k���՘U��X|��v��]���uɷ�q�ΎDX�����c�:ૌ0�ԆkT�N7e&�|xśMaޣ�J���v�9:��XMi��i�s�;��h�@h!ڹ\�hp^&U�52Q�� �$q������t0���A->��׾k2I
Ұb�ZC�M�pQXI7�Я�3�K'�n-1�|zS��N��h=u؞dyh������
�,���#paVO���<��W�^2�b���%�Q8y�~�������Q7xP|I��;��~L#�Fx+O-���rf���s�5)z�Ě�㴄�aFn�Ph�����4XnX\6��E5�BJ�|0�]�褙�,Y��Rq~�%���Nq�+p�r�2�ږ]�/&��)dtw��'�.*t3D�с�}؂��l��E��Jh[�*�<�f��8�o��@����|�BsA(�q��+�u' �3ǥ�*�.�zp|�<~Cb�f��Ӈ wBȏ�΁�'�����9;����W�q-pdQ=�cZ�b�Jq�Z�Pc�6O޵��Q\u?|��ږ�P֪S�)�^A0,Kïͬ�Z���6l���
^~�C��ӿF*>Ncϓ������h�~�T�,�URo^.&ꩈ_0
�t<��C�|��ӟ& 5�#m��l�$\�zl��X��R��_���rg�X�û�w�#VH�D���-Ac�Q���[��Q��������W2�{_Bh�3#/p�b�V��U�@Pe�P-A/���Тy�^m|��Dɝ���E��DR(�w�:�&��	-�x�Q��n��#يC���`�ߝ��"s"��Z�Ǌ�l�1@<T��{�:�9ǵY���%� |.���5`�"����VZ�o[��zm��N����P�п�h\�T��q�bt^�y��Q�?B�KR��g!5j`���/��1"Fh�,Ӳ�oOq�V� հ�'׫���/s�?�P0��g�Z���{�3���D��G���`>d*G���6��}z�iѧpdpI��nQ'T��Sy��
7ogR\���k��~w�G��d<8�����tn�������>2���o�ʀΊ�������Mw|�\��ub\�ׯ�s�k���d}8��O�	���n�k�������ͽ��3�=��+���������%�	��5-a(Vfp�g[j�U��c]^^��_��	���^5�D-H�Ay�qv��R�ED�
(d����+
zi�������
V|P�v��B"�cݖI
r�;�G�"C��t)[����(���#����V�5,ω�� ���tY�z`�=$G�F�o�&���&�͸�&߁��҅���2������o�!��t�(�#�$�p9�$�*�|����O�ߵ�%V�7M�����R�u�ra��ͪ�@��1.�� �j���nI'�5FE{�b��(��n�� 5�R��u��^���	��;�<�O��$*u��T�ml�Q<��2�1!��C��T��V��ʃVv:ө��
H�9F������i���g\�U���V�R��s稩�8a��� 9~�gfx(���mUި�{�6�S�h�베w<.'�M�pV0�& �MizqN�伕\�e!h��"��hϞ�Ҙ�$Vųs��w��Q�]a��됲��l&�d  ,�n��C��#R��n��Y)�i�y��<���9���AK�]�_̸{�|���5�U��:��j����X(.�ԋQ�Z&k0@�&cj���p[�����ˍ��ď-���t,�s�TFA�7���b��O��k{aw�%'8���6cD�^zZ�"�bw+���n�/�'�|�%���?L�J�9��.C(��L1f�����G1y鮺��`c�<��
P��|�b����	�.r�4�Q�I%0���6?n� 
ςW
>�+�F��|�o���C�;��@1c塙ٝ���e��Sx�]�5,U�**�\��,��sئ16���逯�7vw&k����wW���
��,�)K=� �����8w_ SbDld�f�7��K���Z��S�B}�#WOd'XZl�4%Rȝ&(R�|բxt��j�r�a�c��N1�ɘ�)!���K�^��͟q�!*����eP(_�W�H��#�-�<vu��}�C�Wi�
�\�G��h�3�&�5
��D�X�;���?���e���:ݽ�%��<u�v�����z�-z�� b5������E26��4b�Àz�u�Ep-a����e���8�9������'���GQlE?��"k�=�0EΧ�A�[�񍗵+�����Y,� ݙS��y��{�쳂�@8�ĩ郂[w�-.��L��˸�7y��Ԣ��g�l��R�d��?*�9ٖ�4���(�0w�dg��W�С)>v������J�~�ѤӅ�؎R���i��+�a�g���H���-�����hm�+���rI���W�&d{�tskOCY�e
Oo*�s���B�����su��I�I9;0=f�>�r�0��	���6ɱ-��kAAp�"��z!�Y��t�p�ӵ�h��3g��;	 Kl��4믣�����jQ_	�+�`8��:�6�.���=�+�� B�Sb�*g�W^�S�h�J/~w��Xx�>��K7m/
x���� H�s���0����i4Oʔ�}�J����jn�rbP�[��2�ֲ�6�Y;�إ�'�p�P.��m���j�Q�����P����?�K>��S+���Jܻ#��v��ҴE��xΖ3u��b@5!kn�u�XY#1`|Cf�?jק�$�}:�!�%�MZ��ߣC?�8V5j�榢�K�ayJUPEY�[�� z��ˠ�|����I�⁶eq�����(��g���*�^8YJ�)W����53����{T�/�����ʑ�<Y���Fr)�ۊ$#��#�;<�qS�qȡݺ.�����<��ذ���O6�XԽ�ŔKH��[A%�q|i������h�U��|b�,���"8q��2�q��r~8�'\���^�P1��>?o�=m�mt늚<���9��QKf	����mf\>����o� �߻�gj��UJ�F�Sz��:�@�����+I���`hƣ�B�&��{e�<�~�H__B	2l�W���ʔB9C3�%�P�q5�[���63��U���өP�p�%v��N�P������Ï:�����4W=�-
���8/3��<A�#`լ�m�eJ���t�O�u)�Ih'+�m����+A�}��J	 r��$!`\:��]�.�Z�,����ͥ��G�-p�/�Q�F�	�I`�n.�P{H����kBwW �)Ӗo7����h��̺��bo 2n���=O�$v8>�"ŔU�3�h��,%�W��:3�^s��/S����:�r
Sծ�����ʄ��{EQ"�Ǻ����#)�t����v��!��
���U���,�BߊO��-0����M�S�6w�=���)dE�����!�9V�ʡ�;���f<D�C"��j^�Z��-g����C�~Ӡ� ��k��g�,�(�r����e��湖|��}g���.	�4@(R�qZZbj줄�3/�Z��rI�p'[�����gYN��X�����a����1����\��-�7��z���4�}���U�v˧k����P�l����*�v]Z���[��j�&������{�k�=��3��lpQ�����hȺ����ۛQB�[�v��S�E�H����]�}���7�*!��Z�����d�g��d�,�s_�B4}FH�1��{'
�>��
��Q�2f�Py-�&���ԥ���J,*�2���gГ_nBu$�ΡP	���HS�@�nE��YLoh������ILV a���:�����e˘�p��k�n�IW���{�^���@��	�#�?D�W��o�|8CA�ȯ��q��_j��]F'~��Y��\3v9�5���s{���r�[��py�xǋ�ye�����0F� QF��8����B)�W���_�y٘����{F�;J#C����~w��SS��Y���ז=뼗x�-|7�'Ne�tV�)�����{�4�Ye�{�]+�%���i���+��Ŷ�f����ul�"���SL����qI��T��~[���$+�BQ��ٻSb#��ʏ�X�Yt�qm�n�@cV$��T��w�n�����Q�g�a���>���e��
����A��nc�n�p�)��� �Z�,�f��#N󕍥��x��wd����T�H��c rʵDmLo�C�O_ó����_Bb��3�<L+th�Xx�7��T\3��=J7t<��r+{$&�2��1�0�����K�t�H���X͏pi2�#Qm�o����2׌Ti�g�q#^����a�c}R)˜b2aW��W$��y*X%��4x�tU�S��ú`5M�Tr���1 �L`R&r�OF�/����B���N��N�E�Pc��r5���e�G�}�bsd�^�BF,�z��E��R���#��ב/n�.��<vyOm$�m��E�)���M W����L ����($�5^�%��VWP[v����կDAۏğ!�x�a��R�JZ[:��	��-VWƉEM����	Kc6�,��Cg�R�bطĦ��sr��{-g8nX�N	���Z��Z%~�4��1#��q�^�0Z��
�"����8'���8Up6�F�A%����9Y�Z�A@{�=�������lK��.������ߧ>6��ߣب����9F��Q�q�dV�� X<���1p�;Ҡ��l��މ���K��+��@~��:��:��̨��zf��<d�}z�H
+z�X5�0������ ��.�<,��d�ἐĘ����/:_���/�c���zh�-y��YFQ`����F�dP+�������w-��'V�H����9	����6�{��H���O�kR@��	���c<�_���.7:��6�#k�D�(���5,�<qhgN[9Q �K����qU:yDB��	��t��&`����D��6�S�zMp���$dn��L�FBA֔�Uz;#4��n�n�M ����o��e���������=�^e�7M,�rC�a��N V퇡e�W٥��l����DJ�E���\�͎q�Y1:4��n���Т�2�՚�~�QV�����r���k�?��%��<beCc�I��A�]r�]���Q�Ĵ�Th]V�x��1L^V��f�:Q��$������T;BZy�=we;����3T�:E�[�~�wr��vv�0�C����'��{_0-? �CVji�,�ݙ䢛�Q�����0�x�>Qf��1������6ɰT��J�ޥ�?a;n��,�t�Q=��q/~�M��f��<5��P%�z�e<:���{�Ӿ�H.`�T��p�E]؜�ϟ����'�s��@~_BV���F��~m��AvAD°v �̅�$�TDlE��X�k���j9�M�>�\O�2_�{����\��4�aH.�;+�r3/	�_Rfa
��Se�6�-`���(�f1E�4�����+�E�1�W���ފ��	U�'5B�B{�x�����Lmn>����Pa�뗰@��\���
!O��7�t� ����S�9o���Ɏ�p8}�~1`z��/�>�����ˈĦ_��Ѳ���Ft-
���!&����~�Me����+)�LgZ�	��`���|��j�|���<`�x�|(v(cS�T�!�����㽃���wע7�8N,�ݒ����������c�w�0Dik�r�$���9���%(^�m�"��tI�\sK�ӥu1���p��Ȳ\�Z�ࣴW����3��M� .�7MKj���}���U�xQ�B��?ܻ�-Ȓ��� $�=�N}�����A� ���|[��Ξ��c��s!+��FV�i����<�T�ǚy?����6[ܳ�f�r�]=�ᤞr�I��49;�=3�6I��>  G�\��cR��
j�,��C�mk�h����L���@@3��d7jD�Y���͔%`�48�CU����;�����$�9�oW�)����C�����v�份�1�\w�v��d���9�1���;�M����]�Q�q^�ZCȈϬcK��}�C�Z{��a� @�� b���Qj+�������O���*#GTv3���A1�X�=�;��cw����.a���C�"ߑ_|���7�LE��h����{q���'|�V��|�y�*��(�)��:���D�V޿#d}6�s���8�^1�j�R�~��q�-0�9�{-~� q���0!~�h�#��d�p����TZE��=�DXG~=$���v��E �c�����ki���/m�Cb�l�����W�^6�{oݛ�4 ���������_}.t/�dU�CĐ�rq���9�Kկ	[e��l:�0l^���zȮQ������qs^(q��HѮ�^ч����oUO`(����	 �/�H@ጉ��.�9�[�UO5���[I�D�+Z�!��3V�cU��م�$Zb�״Z��If���1��Z��;�m�3}��Ae��*r��E{.!=�8_O�}��k+�h�n�d �l�'�A�PU�rR��nJ�$��|�<y���y5_�ED��Eu���������`fd��pR�ڈ�-F�$�j�;�����P��������EB�
����g�3��u�3����	���=��Qv�I�#A�l+�C9��	����B�cZ��� >�J
��+��r�*a��4CWw���d�+�8J��zМ�����m�&����49�ݽ99mH^��b������%��Hr���ֱ�,uк8�)�? !=�.3�8�B�q+T_�I���(�-�4�(Ǜ���{h��
re�X%5O�����dyτ/��\r��B�T�7介dO�f's��{�S�/�C0���8�����_˞ev1���K�~���د���������9n���r�%v�ԓ{�>�G�|#���
?w��Hù}U� =[-ƭv�+�l�C�ea�i_��[��7Q��9�3|��ɧ�v��\dkӿ��僺�0�s�>M�zL F��У�����⍡���H!� U��k�ھ!�8d�6�����z���W���Ďq(�s9" {Q���%�l��W:]�	���u�E��aI8�^�G6h;��g���W"�����j^�e��_l��H<W>	a���iP�q׹y�}EtD�Y����Y���^�Xo���
`]O�:���!$�}�L�b��w�����Grb���	,�-8{0�H{�O=��z��CiQk�Ph�~"�W7N���uÙr��7�$?u�x:d�l�����ay��
�b�O�2e*�}]���d�7̺��J�ٷ�R�Y
 eO�����a�5lԯ����F�w��8�{��"[�获��M�ʳ�(�c��3��W�̝��e�`}Ѽ����)�R�Ǝ���dc�x��i`�EB!��s�C �ļ��;X����7:� �ie����;�Q�C/)�B�c�	������q7���EF��-h��Z�c|5%4˛��"�w���-3�l���侗�� ��ydL����(��O�=jh��Z��jb;q�/QI����8���N�2	:/���u#몵�q�T���iv5]K�7�ӯ.J�iF ��Ae(.6;�G-��bM_*�ǻ�c��A1ZQ�)G�Σ
Z7���d�A�=���g�q~�<�.A�a�,>��2 e�¤�ϓz_���D1c�C�5c�a�n�
�w���?FB�'(<@V�(\r�G'%�6<[��f�>#Ӈ������$imj�`y0���*s%"5D��p���q\8�zS�e�6�P�ؕ��ʊn�i�%Fx��D���IM�Î��n�Q0�d~�Y	�5L��5���Hĺ{���Fr�(<ÁhLO��h��-�g|�����mDaؾbo�&�y��U�=�܅��Hh�{������m�j�o�$��{Q�����CĀ�u�����lG1؊�>Q>��;w�nTDS�{��E���ed(FkA��z</'�CL^<X�vZï%:����6����3c������&�����{g@;�[#��^pГp���q��[���eO�����[��o�Z{[<Z���x����Rj~W�mJxg��7wH/��W��\K����tU� ��b!��Y����o��<@ދ�4����L��I���Qq���I)ْ(�$��,!^
�#��J��%�'};xĦ�X/��@�� i��!��?����ў(��#�d�9J�e�E�'gI)�og
�@+�ٽ��B��n<|J�i�A�+t�	�%5	(ū����IZ+��1{����촯����N8����ą�Y�ƽ���Ƀ�;"�c�F��*2�+�i|¤e����o�O����W�X�>o�G��_/�XՔ�a��������6�P��8.�hߤ���Z�:���R�xy��9`�P֜V����&!	A�a�n���Xo�8�%��Eذl(V6k+o��û�a� �%t�I��.�K�4��l��Bn�\��{wa#[e�C+���E�Yg{.bG��r����#�{�X�x�g��<�Q��2�!*G`�WY-��:�s[����DAL!{���������\C��N�6�!��ΘWF�#'�:?���IZ��$8���Q+�[ֿ����6��\a.�vD�����
a̓Ty�*�h�yĜN)���	�K^��+���ؒu�H&�2��d�ڶ�Ԗ���yr]��n���K�3̟��;��f��D;����B�����\_�����-���0$��O�c��OC|XNGlp#^4/�[HM|�@-�ê}�X�#���!Oo��(� *�g�|C[s��k!�^�>���Z��Zt���0)���%�2�g�O,2]���vj���oN�јn�a���� A��63y�0pv��h�/L�n��Q���o�6w=m/g�Xvհ5��ӫ\��R뱑�tǳE�
}�T8'fL˴�����\}����,6�y�3K��ʇA����I<Aq �w`?�!���5]f�:_t��[���{�*�0�.��$1�c��x�?��/b�_K�ZY���D+,aObH��K�k���ݰN�zc��:m@J�%~Z���~ %����p��?Ϋ��P72U�gZ)V����}'b�U8DH}�]�sr���ڇ�j&ĳJ���Y�W�T]�̔��+�P�]u�v�8�9�Rl���H9����Z.�c�]��a���#����&��=��#���D˅!cw��;հ����]T��L������w����= ����r�
7�oϓj�J7ڋ>eJ5d�
����5Yr��yt)��ť�Ǯ���1�
�_�d�9�V��,R���G������C�&[�B�)\���u�7�?���I[*��㌴�s��6e+��W��!:O H��"�ݵ�,0຤m�����k�>;I��r�,��=(��@�W$�.S�$%��0ޛ�K����/%�J8f�������t١AW}z����Ovx:A��M6X�O-��\�C����������dh[���ޕ>&2�:(Q���Ke`:�Tz+.�#^ϟY����>}_"�IR��Ć+Q��K�K�M:���qH}�=f��3�lS����bcST�����hT��s8�ّ�>�3�����H�(�lI���������[�`���vi�����,ꦭŗeP/6l%�G�e?" �-��_��x�Ĵj��%�X7wF"���SDז��r��̇JĬ�I-&�)�;�Y�t�����=�#����NpZ6x�"�L�7�Bq;{��i��o*:֛N�J�~ul�#IAK�a��_ɿ��#�95�jN�ʞ����.���p@�y�`����D�����]���C�l�\�c ٭"�~9�G����+����O�8v{Pv(���gL���O��JV�%U�\�{�
�bc�Ɨ��
+�~ֈ�5C z���h�F�Ҏ��Fj!u3'�� �>	��WkIN�d�\^s-\�~�F��W���� #���i�Qe��v<״�.��V3I�bv�aJz�{GC�[ໜ�>8���fu֩�'���)�S��`��4�����K�3ҳY$�i���GC����X��@uc}7k�s��ӆ�����W�]E�$6�$O��yރ�CfQSL����=�5��."n�poF��@x���ZA*q&�<�+r6j��S�I�ڕ��ؘ��,������=����@gJxP|����,z*��ߣd�HR��(%��T,�h?�E���W9O�ղ6�|�������㹵&r�UU=��,�"!���T��/F�ճj�7c�ܧXe����(�$O�Z��%a��>>�mnq^8��N�`�G\1�8�@��D����|�'��Uh,�h�(��ꦕǾ��9��[y�A�BíbƷ�w��#NWu[L�tE�ſ�X����[�g�e��	�k�5p��)���-�/�W}�69�i��Ж"'���H5����v1	8��I)G��[ɟ�2��^�G���:l.�������R'������ �h���k~����pp�oB�Rz��D�	9�
���8zmX{2�U�����Yf����^̦NQ\�O��1���)�񥽡�T�WO�� ]_�Z��v��dD��¾�������UII�Z�}���_���>�5#��&u�/�'�L�@����D����iK[�.�<Xjw!�A�tjfEi�g�����[#l�ߩ�V����1�^܀T"�r\lL��<1�܃_�j��й�[簅�a�[��/i�k���W:E� ��[r�y�f�e.���SU�~�HE��!���s@*�?D�ޏz�d�<���y���>�넔��w�"� H�A� ����w�7�4��!*�n�3�9aPPgO[�Ш�1s��2���Υt�+��]sBܞB#��Qh��´��|��l��g�0G��k�(�����C�	�곢hi\����Ô3}�&䥌���j9I�E��3iH��K�TJ����݇�Th�bR3�������H~�B����;�PG%�ԳGپA<���)E�Z�-�h��`��
��=\-���M�WF�<�ju�P�Ŭ:���e�0��{�l\�|[yR��l-ǟ'��.eb��c��S?>�� �<�9�8�=ܱ菏�q�İ�Z���v5������gp"4�����ȖS���0|�����4�0�wa?ms�Y�����HChA(�frDZ���,��9��vv_�m��k�{��*������I�<��ߜ����O�iXS�CXM�G�'/ ��PJu�"ZKd����.�U�7xWh�*��^���|�~�!\�|X~"��d%�B��~��x�Yb�_���ze�/���yU�� #��P8�=�#��A1�"�};3��ϒ�y��TP��Ծ�6�̾8�U��R�*z��6}��-M���ՀKxW�̣ô̫��YN���w��1 �K4:�L d� ���|���L�K~Gv�푬U���ps:b��}��@e�D����,��W�m�`GVD ?����/Q++��Y���Ea>��egH ����nt��N$H��Fh���#!�#���.؊�\� iG=�Gg�B2O[��6���OE(��i5�*ơ�",We�{'����Mi�U%�����e�D���	7�3JKL��s|m�z����uZ�t�5���\���95g�@1�!yQv[�a\1ޛ,�tƖڽ ��ܓ�V�H�BBm$nCB"��:l1�n��$Ծ����a��xT�4���sMPcso!ԧc����rl�خ����Zj�%�4��e��e�É*"�/M�T�`u�z������6%�E�H��XP�my<�B�X��9TT�h��xF������0��̽�w��+�V�3�ل�W+P�L��E|�tb��uG�8/^v��10�w���U��e�Ԙ�{KL���+�X�X�#|j&��@���zf�O7gq��NvC�n̈�Y]c\.I�Ġ�,���n�ċFa�����a�~33���>`��\�m�t���?F
њ)$=���S�Rm(���T��e�[(d����>�xN{P��W/aH�c�!�����������-]/�Ȯz�����@n�0�����ɚ�U�kb�J�C�+G<_�\bI;O�8ܗ��w��wI�����p1��z�&�R��a�ԋ4і+Nt�?<�c.S��_G�^K�o����_�KS裳��%Z����k?R7��{(�	��u����[Z�J�S���Ss�l�Q ���Q�Q"��Ȅ1YB_�I��1�l�Uf�5ͧ��S�� �B�ʮl]<�؝Xw��+�Y[1@_ �B-������Qt���㷡<��-�H�P��>�����Y�Y��|��N��m��
�s� ̓����M�E�8�&���`y�S�MMP��*�iXf�t�Ġ�y(�	�:3{Dq܃������dXi#��K�o�]m�8y�� 'Rp�\F_��(���$��x+��:t�E{s�rZ�"xZ��� gʖb�g�9=��>�A�(/�˾N��A����������̾K�4\������ޅ��L������͝Ǫ�UN������5�Vu�����:)�k·���4;��uF�}�[]j�i#����� ��I'�$cqI��O�C����틋Ijv�W���!V6 �zQ��Ϸ�Vՠ2�����e�
�4�H@p|���Cк�ڃLgFLޚ)T��6m�1��Ff��o7	�+I� (�L92A��6l�E$�n�ol�N;�K��H\�!��}z���$[���{r�n�J�K훵x�J]��l���h�+���U�uN�]��\�ǒ�zOI��8��
�Bg;׉-#z���rq��N��(u��`�A`e{�p�K7�H"�^L�yE����*����*� �����E���I!������Wx���|E�mm~���79jהk�6"ڻ��� V���4��^�ڎj&s�[ۙ�k��ȓ[�˨�!�/�%�>2BÓ�X���H$�N W;��L�{���H����~�!���U��b��Ar^��c�'�<�,���¢�P=Z�+9�b�j��BǑ���]��ƌ���VOׇ8� ��3G�}N�~/-�b��o��B�;��ߚ�'�og�I�;���M�l:B�p�2Gp?�/���{H���B�&�!}&�N-�J�2����tZ$�N:�7nK��s�+���D��<�
���3`XaA��Fn�>#ɒ���8�}�Cq٫y��d%��M�[S���4�}�+� �����"f/� l
��-�H��Ӧ)g�PBy�f/���:]�_0���/�a&�pMbҭ笑�ho�8I�<qE����z5���b�XS�]_����lܤ�'jA�q�V�!��m����680��К��yN��@�mw��)�1�1f?ٓ�$lvY���4-U�+Ҷ����S�Ҍ���ʞ�WH���d�i"L$t5H��8,T�NχF���7R����zHR6Pz��u��@�m�J2��Ucf����g�~������i�O��k>���Y��)G�:�b��Q�mR�SaS��+bIP���zyb�L-Ӓ	j��Ǽ�0�ɜ�UU��QQqt�r;�"�� ��n�}~���x#����z��dm���9�9��֗��b$�H��E
e��%��%؊�\���.[fe�HM&��z����$$?�2��0�^��1@>8�1 ywc�c��9XM�@L�n�����^&��:^눷��oF��w'��^ ������OE�rJ%��w�A0ES�S�\�)�F��$/���V>�Ut�7����sN�{ �X�F�.p�Z9������iW������'��t���-������}��pSny�ʗ"L��}����|�9�\j�O�
8pH�x�ji[M���xW�az �ޫ�],I�Hb<�
���uU�q��c��I�PB�7�//�w:b9C�⌖����f\�G�M;+y��*����ˈ�j�N���1��K�/�g��U�����K:a�ԯ$����K"SU���X^[�M�8�7F��Y���-1���A)�8���&T �x4�cY|�5�4ױ�N�(�ԇ���'W�n��f;���?zxbJ0�- wЄ��o���7F�&�����;���Р��o�qOKt�}������C��N��
HH�S�EW}�r�j�QQ��c�����_�{��eR�8�����Dqс��-�,+��j��R�V����1^��z��m}�=)'�����%�����F��s
\�dH�j���%��\�kU법�L.b`sHlK}^x�.C��c��i���U� K��� zk웡m8��[56��{>k�Z�"!3��Vtҋ���vڮ���3B���?��T_�
+\'�Nh//_քح�8��II�sRD��h�������2-Z�����X��vkD+���7˼�=) i��/��J5�ٌ3�'%!��A��g�n+WBW[�I�:R8w�_-�Jf��c��g2�X.s��Z.���7�y��?�.^�{�����������'\��vQ!�E ӻ�"ů.�������Z�4?���ц��%�C�"��фI��Ҕ���،�n��`6�����F$���^��=6E�E>I��TV���p�+o"T���D�U���4_���z���RRb�b�W����sƅr�s�͛��7?������]��V��̣�w)o���7Ӌ���	�!-ߤ�?�ћ8�qڶ���Eͧ⢿���ib�����J�	���*�wO,�eV�����_��^$��5z��f+�� �ѱ��������t��!��ܺ�.� ������L�k?�0D���Mz��\�酲�^�3�~7rU���{�:L�E�,&�������%B-L���{ ڭ�;&�k�#u$R�$��R&�����+��Y�c=�_�-�Q�T���P)��#�g6ɕ+����ן��5>\�a�ě�t��1���s"����T#�9=P]�Omâ9�g�&[%��~��4V�otxA�Le���\1��иB4�e
4�P�?j��b^��M��vFM�E�+���e.a�E��9���CT���#��܉�TbTB�*swVe������=aK�J�3�Э+�&%��%���Q�����+h��e��5Or�����E�%�	����y>]/N��}�T�����'��/2�P(�N�:�L�S��PE@v~�4�#�9W(�$���=z׶_�C�fkx�*��r��+{h[~d��V�L.\g<�
ԡ����f����{M�v� ���`�`S��=Ynm��q����r*p�_L���pS� ��Vˤ(-*74���֠�iu�!���ل^n��^sS+O��j�+K�ky��bC ��0����#%m��ጜI��UH\�d�m+Lgg k9jD�1L�t�B/!�sF)1��u� �{C��<y!����9l"]��~����]r�����ᚯ*��χq;�	��V���R9�b��v���mW����IA��uH��u�%�ߋ����Y��Ζ@+f�c������`�TS;J}{��$?Z[d ��"m�9H_�3~i������<�`��P� ��!��$&.j�DW9�p,��OH�����|r��3c�ݐ��x�}6lF~��Ó�]`Q1���%�~]��s�>B^ ��71���o=��ϧR/�+����@&��2N�9SA�\����7����"Xe])��_o�nGt;7cg��F7��\�Uw��'���|wĻ�P=��6AK�6��<�j~�>�:�ګ��i������f�F��HltE�wLb('a)�B���q��
�@,y����Nz�qE��&+�Z�\S���-�c>�#�s�U���s�	'>@#z.�*���0�-�b����-|V�Ƅy��N�7e�ַ Z�w��.�ؽ�$�,�pJFLc_e:��	4�۞�4���f��ߦ�	x�i'(�ߤ��h5lH������G��9	�������#=)b-*�J$?���z�a`��.˂ad�K�K�]c���}���DB�7�G�x��Cr�T�<�f��՝�f�BUL��.Ʈ�p��1#��E��ZU�3�+��E���*R����С��DKN�,�2�Ub��ԚO�Q�ֿT8!�Dl��k��n��T�N~;�w:��,Sk6�4���j��f�{PM�.�:�╇�A�����������+o��-�?�t�����B{�X���Xi��%�+�%����;��(���'JƱ���opW�2��^�<n��8fA�~}x���sc���ϭ6~l���Ĉ	C��ؽm�d�;������i,N�G�nS��<��[-,������>��i^W���,�un�ۦ>�
��GY8�|�W�L0#JJ.|6xs�^4����� ��Fzٷ���FC�#��Ra�s��v� ����i�����HD<�'q�*&�����YP��_����"��x�U_䋶.R�&��і9�lh�h���5��.s�݆���K�yի�#��e8"{s��&��^�"�ç��'��F��h��}���*��SY^G��'ঞc���� M�ZP�t�y1��7O�������F`��D�Yf���K�~��n��q2�����!0})&�fc� ���4���6��P���Cx5ϒ�+�F�h��� I��%��Z/��L��!u��e��b\0eT����Gi��r� ��kH��k�;��?����c8���m�M.��'P
��x�F��9H�Iю�-B嶼6������	�q����hy�}���]���R�l��R	 �u�,g'd�S��`�՞���@���@1!�?�~��%��N�-a��qIc[Faq�b��X.�T�(���	��~ú)��%�&��ޯ�����o�:�:,�T����|��]���oa�����b��Y`g���@b�؋��PԤ���V�k�ݷ�l���7f4,㘵(׎AI�b^�@Kj���y���Ҳ�tY=�ŀ,b�V�!�&ޙ�:�c���JV���#{�^ך��@昇<��9ջ�j�#ι�;@��[���	��jL2��:V׈�uÓ�;1:�m8�X3�ͥK��Y�o͹�m
�*�0M�� D�v
��n<��Ќci���F�:
<\��J�yh�ڍ�����v.V�d�z#Ԫ�o�<� =�uX�J/<�dL? O���F�����,^=U�r`h��� �Ro�t֦/Ɂ$f �*¦s��?���������|�%���F���2�z������E	�m��!�ot^�ȱ���bk���v
�(!G���A�o������9��}�l��]3<��F9���[dՙ���(�����1��f�U�X��z5e���Z���EP>H}o�:�+�n�e#W%&W+J�6��&�|���t�a��"�٨R`�r���ݦ��I�֫ŀ�6���~���A���/*Q�ۄ�u�:��^����~8$Xzk�39��Cla�O�2dW=�mn�1�n�.z�uaFM�
��(9�Ke4��؎�k͉�D�[5B���%�~7L��~�\�/��xNջ'b��/j�x9/�AR�r�����y�M/ry#�it!.*��R�Z�m���~c���Vz����?2�{�ڄ	泜�t(H�6-_(�OMyF��E��d�X�&X6u+���K��h)�O2lsί��P^Y�T�Q��xi7��*���]��<ruJ��D�N:�@�	J�g����:�����|�^O��TV��@R]�Z0�$+jI��v�:1cv��ma�4���x"ev��I$ȝf�k��u2B�j���	*CE��5q�q頚@,1h�.�
c��A�)!Ff%�����������?���$}�R��U��[�� Bg�\�;m�IP��V�zO�܄R�{/$��˶��!���.8-��"�B~��_�;0��{>jDq� �9O�y5|7�����ΤR�W���k��G�z�Pz#�C��ڑo���KɊ��cq��n�Q�6�A�� zY��X��Y)�������M)�@����,w�2j���9�%{9r���b�
v
��x�b� F4�i��Jm������M�h����	w��sԠ��EI�ҫ����)7Y C�.�%�]������Vo�����uO9[����l,2`UaKh;p��,�V��_�&���Ƃ�E��-�[)�������)�r���&��d�:Kgˤ����!���d/:z�b��F遡�1�1�?#-�z���p3ٲ��!�zlr7���2I�/�uHjP/���'֗ �9�s�΂j2�z��jU�a5�z�-�W�+*��y�G@p�<��JH��I�\�k�c��~��	-����.����_/m��g�wj88"D�F�L�{�%
��U����ݴ_���ô�j���V	v�!�<tء�&ﺳ��Mu���2G؜x�%,�j�a���_&����lѢ��__nAz<�s֩{�?O�4�*b�ͼ�ܔGR}��Y���Ou���ϳ%�C��+tKe�b��E@�E��\L�����^�( ��yܔ��&�����gI�dEz�#W�I�$������{>DyV5JO����H���~��n�S�o^_����-�".c�·�Oz}p�T�L�>1��Eb���x���F#���D��
6Bi�gbr͚�&�Q�S뫙{4��<���ru��,>yl���H �x��)�����jz������-^/� a���>��Xe�-��>S/Vi6Gr�=�; O��Q�N(�z̮�F�l�	�?o�ЦRA����L��Ga"M�;
�+S)A\k-t��c�b�|�>�L%k�Oʊ�Y�6+��	�[�"�3�G�:q�h��w�ֹ�!3��2E=��w	���	�ō{!Z�'����W��5_�(U��ͽ�e���ʄ����R���ObQ�I� X(�j3>J�dm#�vUù��TWz$| �e��R_&=�5�Ss��_��뗸�cA�L��n4.�U��=5\7!!�I-+`�t�^Z�{����O��f�9�����(��T|���q��uD�|?�l�@�^�e�ғ�2;����r6Z���ikiq��F����sTd_���� ���r�Z�:��v��i��w��K�`F���P��wT�� ����^��vF�Pa������rm���RL]| 7BQ�y����:<Q^?�yR/{�@ې�j�?R'uq������:��8KK6W��v�S7<|E.\x�:@,5��0(�?n��~o	:��̽v��G��S���.CtD&�dy9��;I1�|�%���{O�a��_�����L�${z������k�t���Z#FD�L��q9�Y����L��l@`�D����{��aU�W�o[n��hbP�~JR����Ľ������[/gQؘ��{���Iyl#A��	C�Iqz C�T,���[5F�U
�|����w�d�d7��Ng�=mI]�s�c�K��ǉ2<�acށ���m�P�4[9���#1�r��s<[

I�)h	芬��q�v�{���_Kz�u}&oL�7��^d�����o���r�?����+ʰX�?(��bhnfY�A>�o��|h��+Y��-�A�ϓ <s酬�!���Nb��e�d�k�\D�:�a_Jc��yŪ�f��I�;�qi����{�q<wƹJ���o\&oKKI���'>;d(��Wx1(ěf�x����ӆ�ݚ�3��5q�X��.(�k���4f8�#8{��zU�Q�?��Q��
3Y�D�=�N�A3Hh��%Vs�P�e]�y�����
�(^��|Z*�xY/�=�̎���_�|m�)g��~���mEVEjW�dL"�����W6�����R�>�#�k��[�`��͑4NO0���߃��>��I�)syp�#���Z�{h�/L�:*D���VF�6�L��m��`$�'>�;�;����)|\��[�z��p$�b\D����<�lAP=��r"s��ΐd Xwt/^ہ�J<1��
�>���:�=���J�_���N�+�ih�:�L���C�4,r� );.�%��l�|�� Ԙ�,��L�����Uo�!�;��~e�3 �;�B��w��`O���#���kp`����������mf�y�]&��7��m�n��^9'�i��m�{��3(�s%3�2��	�E!��-L坶�&�7�1�
`��Ս��aY��z��ߧ�}�w���:�� eD��ک�+�%W'�ee�}`�8���� ���fjP
{�5,�">�R���^_�M�����W#�����6_��~,����|��D� ��h�v����%,��ԯ��P����qz��O&�V b ��r���#So����+ܠ��@�0���F!�y���noK�;[��׽���<RY�2���go�'M�F�)P��7S�o|j�E~GK�ˬ 1e���Sʘxgّ��h*J�������n�<h̊a{�9����I�p�GH������d(��E�x �%r�j�ӹ��S�*����^�����8�����++A�$浕|d�wY�Fd���=m�_���f:gZ@g�2��^#[%<���QeDmC��$��|��$���¦���@�1J�u�\�	�9^j
�#@��O.2���}�߇U����8f�?�l��'e�a����3����/�a����Ѥ�(�)�?�!8������5t#b���lB�՜��;
�vMW�R�����ԧ�cB������!%5��K	����p�.����S7s~���/j��=GD�U�=����W�}_e�f��� (��t?�GV���)�4�
��0���҂g��u�6L���ژ�o�����C`�8ڟ�J涡�Z@���p8Łi��Vkud�H���w�"@1�"��ϯ�{��{"�T���2�WA�@��X�j��I��0�	z(� ��$�So2;C_��.�۬E�^�U��8�Kc_�]���z���������5�m��G��r��YND7��9�}nl|���[ÖRU�[��-Z �Ta1�լ�-��cq�S��ۄ���G�7C�#h���A��:g�P;�_�[Y�����ZW3ٿe��&��Q �Е������KG�������{�~�c�K�� �����2if=j$�N���ـAq j�S��( �#.,��Z�)cgN.q�hriH�����9�,�z5�`��*�<����B(P	�YNY���m���8q���u���+�<!v�'D��?�r�$�СT��=��մ������z�m�9dj�љ���*h�MoS���'�[�������_�>Kc��#�[���BlU�6Fkzi�&�Fx������f�*���*r���N�Q����],�ŝP���F'`'��=�1�[g���ބY�QF��K��tCq�r@u]c�Eo��-	����s-���)���y�ų��$�2�`l��t���A���>[y��(��͌B�s��޸����d<XO�"(��2%O�z��%��n�g�}n����9��A2S ���E��Þ��3�="�3�����f�8Oe�`�%��[�:^�	���l��Nr���_�Y��C��u�P��_�������<�L����ZxBѫ�:+�R��_)��$m>$�� [��FVJ�k%|���DV�]\t$���>L�.�be]�x�jr����yK肬;�Ֆ�C-���~{�O�pr�u��9"�Y�}�U�P���d
Ol���_J��Ҳ	M�<j�l�ē[Jm�ESV�F��7���
S���I$*r�=������y͊��Ni�4�=\��JCb��g�ƺO9dvH��H�� #����f�ҐocBj�0T-
IP�A����&I���X�v��{c�3���$�dP���q ��@�w�bP��w�'Re�Iz�r��<)Aې��.�����<��K�~���U�'��JO�/`	��!ϙ��9�e��V��+�C ��Vf���fe��C�t6$��Yse�A'2����g"Ƈ���H`,�Tϫ �S��}���C�{׾̀���Ja[P��}9W��8����ߦ˗9������/g���n�>���ٌ���6D�OY��������Py���,z�^�/�����ϖ rC�L���|�)�ǎ�fH� X�B[��IF�^��>�o�����
L�u��b"{p���@�rNZ���B���k12�w,E�q��ϒ��k��t�8lP��-�:��#VݝL�ei"9y��W;�'��U�^��dw� �Ul��T������%�X�a��VF\~|�.XAZ�Q؊&��^�Ir�s��mNI�A�w,��=��\籯Cp�tn��� ����bSY/��4�㺗d�4��y���^?������oY�z��I��3ay ����,���F���,jj��(-�s�<��n�`�E�F!�t�5�Dh���
�-Y\E�p��$��'�}�ؐl�_�Մ$0X֐x��(*��;����*�$*G�L�g�{q��L��zGzU���s��>�$8��C �e6�Ys�au}7��?�����A�Ǝ�ʈ�؉�^h%� �֦"Z���+��l�K ��������w~�<���\�I����I���82�׺�ui|���A�:)
Y�|��}�SQ�AN&��b�7?%"b���Z�V�"خUɏ�;=�3��u�4��ɫNU�C�����1����oʆ�4#=r�a�U|�����<G�iڜ�B,��?6�	5�����M���������AE�#�
�a8��H_��֨����JS����u��ڜ�5t�y���e�um�{�Wƞ�n5�B�}l��K0�b������q��\�w�[��<��<�Â�q:��Kj�3��)p@�>*	���'w�(���ٚ�����:u�fY�@�<�
�~�g*|JT=�a��w��C�E�*��Ot�5+q�4� �'5����M ]��G^	��	�b����u������?��0}�l=�緰�e��M��nY��%����$l���w���DN+ ��s�p�=�i�>A�K��4J\g}S�����=/��>~@�Ju|�S��1o�ү� ���!�����4g�gC�o�!���[�3$K��PW^���Q�!u�Z���t|-J��x�p�[�(���z�y��!��ш����W�8��~�U����F�;	�'aYeSO��q�SPLgl,�jA���m���糝Q�\�t
!�
�~t��ꪪãU���6u�	H'�'�1�%�km�m~=_���f�o���O�Z�P̩Q� �9�1����T����ה~�`Z?���hv��X_3�d�'~ �M�el�HT�`3}�}�Y/����h�$���*���'��
f���������m���П�?7Y�l �&���� ,Q�q����R��~�qР��2�
��(fr�I�4%ve����&<�Z�c*�$��VF��`P�T�u����k�T�YH�0��{Lޱ�q�?,��N�4݁�l']\�[�"�׽����3�����*���H����Q�17������� �F���Vɦ/B�����e�z���B���ɃAl׌l���~ٶ�9�$�Hܶ
i��0K�_��/�	usH3D�]"~+�F��o�z�.k
`��_L���4+5l�Т��qK�M�`ϩA��Bga�J@�Ds�ר5
$z�N���
���)_� �j�{��h�%YKvH������ʎ��8K8�ZL�:,������^(V���M���� Ă�&k�� )�\�[U��,�6�J�(�l�"�:�P�</�l�	Y��e^o,�5�&{I��+BL��a�?�{/�`ʠ�"�`��_�{o��lT{l×b�[?uݳ7�H6L�癩� ĸẕ�.c�C{��9���3&��%'��x/:ߵ:�Gֵ�$);����~��J���?H�J|''��D�ח �ዓ�LR�D%ې}��V,�-�:�P�xsP�F���ۘ�
�/��橔���a1/{	����/�� �w���3�C�ID�G��6Og�\��e(��f�}t���0P�1�O��q��'�ܱ�d��n�'@��`F���R�ۄ�H�9�����k�v�^�A"3�+��ү���S��D��U�⻺w���'�H�իz���R�A����3n�J��	|O��=&�U��OΆ?3/(ՔÀ<A�u�q�Tߠ$�A)=�y}G:DL��{�˴2�7� [�.nX�p���>���Oo�nP��x�v���bF}+���=�EGXr�:8�����	���'g���3�'���q|[L��X��@��,[��Ik����QN�x������@�f��r<ﳆd�Wu�2@�A�$�"�M�5�����������tg�%}:�9sy�h�V��a�rΘE���Y�����K c@�.�Vo�!�3i��b9�ٙ����]���;=Y��҇덣��G���5pu�L�E���B�Sې�����'|Q��Q~Ll��O�Q��F�$wm�r��Nᘨ�jJ"e�I
i���ml��/өZ����Q�vI��[�	ƒ��l�^������aW)'F�}����g�~.��?��������i��M�S��A�m~K��\n��J#g2��6;����F�	pHc���</8چٟ��_�����V~��\Z�l��Êȴ;.���r���'��
�D������K0a7:Ԙ1^�!5#sj�]�Ljy`=�,k�_	���)�dWZ@M�"�>4�,>���G.0}j N  +d�~-�`���SgM������	�mr�c(҂�ZI[]�,OP���tӴ��m�ഠ��ހ�v�^f���M�p��6z9(C�^o�Dt�N�gi���$<��LT�j���"�L��.	�n:Ctu�P�C�x@g��U6� �\0��TA��| )����w�m���s(��U�S�!@�l�mR�i0�M>�UOEcK���=<���L�`��K�6�ɆeXjP`G�{  떥.TL���FVvulòK��?F��,B/��`�%M�=~ʵ��ES��P?�Be�F���[���Vӄ�Ujr�h1+�;
CPQ�%�<}Y-�bkPJއ�IQ������w��̷	ƣw���4�(R�M�B-}Gؔ�#��%��v��}4�}Fc�ġ_i��{&�}IȢu��+$��B��,!fW�EjB��.�HL�(}p
hPsM�~md�zR����_o���IR"]���5��e����Q'���(љ�MKv�M���ݪ0n��6)�����/+*j�o̊�U��D6X$]�Ak6�ͺ���z
��D�W5�E�V�28�/*�Ҙp�%u�O����t�}Eđ����T:
���7�"~XRJ<)"W[}g�xb�����i�W[G@E�o��a4�t��;c�o��n.!�sy�`�0PެK�!�{}Be�$�t�%�j]~��
��� �cu�[&�ʁ�5���"�̔�E�w?LԒ�N��r��g`[R��8�m�g�ߝWŬ�)~��Q�fݴ�JlI���_�pJ8�>>���j;�)D�����(�c�]�6�#hp*�6Y��4�^�e�n���Z�ԡe`J��+�HVr�����;1c;�Yg|��Ҍ�i����o��Q[I����.1��ܜ7ϻh�(+YUn�i�7�>>wa>��đ�St-����)}�B�7��J��0.u���_�g/�&�j�:��.2&�'��=�i�q�
A�d��&8D�7�!�nXKz�]H��I�����^�EsN��^
��R$��2�gҩ�vT9�uQ�mS)"N��]/�_KKp|#r�H�\{�$���y��=��.$We���;ɼrڡ��/���}�_?��O'K���d�	}tQ0*�'�ͻ�`��Jţ]��F�2l���+,+����?;�A��?L�:P�c��Ō���X��UH4U�&�0C�ytR��3V���>�jU�߫U/�
^��F��a�\���$rMQ���$Ҿ�th�*�.�F�r���Y�}� �0���#H
:R�� ���x�a�Qyg���B���=�j/���0�/���J#b���ے�?����r˼8G��g]��̻�rO/!��]��`	��术�����uM���^�ОG�{s��p\�|�.9*�1��N2j�n���5M��B���%P��&Ӱ�δ'6^�&y×n�6��\�;ҭy���)>�����X�5$�dӜe�3i)��#��W�����oz�u��7&Xе�As-��<�ǋIG)�'t*�[�ȼ���n�8��U��v�JS��.5�}�x���E$��0�48U�D�c�e`�5h@�$~�������ǀa��fB����h�ݣ��O��1�B"�U��>v����ةAyNE�t��	��j"<7�Y2؟1����0��[�@ڋ�>�	�G�_���)�����G���k�����{���Αh�/���@)�M������7�w�s����o]��+��R�\�	�.B]�݃9�E��𱐴�����TfT0��m����T�Kj��]�Y֭��R:F����3�<�^�����&.�՜qDA͋��yH��pg!' ַdi�7�ݛ��[�´Ҧᩊ�D>B�H5q�� �h�$.JX]��|0��];��MO�^]s����"�\`)��L��>p1>�2��HT�4:�H�wc
ǚ�y�J,�h���n�9� ݟI�dE�8�-�-QW��nۄ�/�<'��Vꇕ���B�M;���e��х6!G{�ϙ�-Ϥ�mU��^E#�0���Ɓ��;T6Ӿ��H�@M���f��a)Q Е��Ɯ?Q��&�eCy���`��f5^��
� �HB7���elE��ڕ�:#�H(���n��yV���b�6�X�o��,��,	ߑ�}�F����p��(�~e}{7b`��_��B��U�����a=�;�(SS�L�ah4����2z�ʗ�)��Q�+��A`�~��j\��d�_׃J�*���ǆ��� ^;��&W����&ϑ�l^�N"��|W�17Kg����/0�ؕ�����fb4/U:̎��ߎ�g냗 [c�IxU9m�ZmR��>t�c�3�?�sx���ڝ �ٙ>wW[~Z�
�"L��s$Ͼ#�k�YG��ơ�贐˥��l����X��0��R���VM�����S�YS/��MɄXIV�
C~�Т�)Z��W�ԩ�ۆz��c|��|3'F�V�Svk{D|�%�xr�ѫ�B��"w�R���di�wV���?�஑,���ԣY�>d��Z5;��Ds���̀��O�z��6���'}O�3�v�Hq���CD�,.k}��⫩�Cq>���^�M����&�տi1_�\����	5:��Gr��C�(	�t%(�������u@yC�vDf�u���R+S�H�J�X�%�q<4����\-�Bf!�f��Z�P�u��\qb{T0J�C�G�Q�G=����`��ο^Ol��Ŭ�Ӹ��{6Z8�G��&}��.��=ZG�)svJ��W+���k�ϻU]S���{�v=?�t��EW��^�:з�D_�iT'L[C@�鷀�
�|%t[컁A=9�<T�Z4v���"-M���ˬ�Z?��{_
M|�����R+��#������ƛxU�tp#�ٲ�{h�γ�Cf����8�Ut�����jj�k"��(a+,�Sl_�O�z��<#T��R~�~8u*ڼ���~�Lx ��C�8�2"�wǪD����f�7�Z��W����&U��ݻ�n��FN��/TW��S�䉳��#��_��C��~J��T�abw��3�N�E�H��i8?6�u�5����t(r�&q�%ܩ0��)�^�������˙����Kx�������S��d��5s�����?a�xJ���r]w�j7Vq[l���,E̎�ۻ����Y���&j�׋q�o�!��5'���a�ĩR	$:v�ciʾ��T�M!g}&�W�?1� �"�F&�U��U#'���r��c;]0L�J&:����e!�/�t=�$�{���kv}F7>�=p!�13�����^a���f��nm<������_��\���,��V�u�S��QW�Ù����pd���K����Ϩn��t��_�'�9�� ���Q��c����W�����i�l�h�>��pF'��G[D�G����B++�'���Z��d$ue��/ÇB(!�g���0��;Z���� �ߒ�������+�V��_d��~2H��X��f�ꇟ	pr����ѝ6�`��4@�_�&��Be��")p5Nq@lz�O!s;P�W�h��?��-n��Ek���Pkh`R��CU7�������(�F�Y1�tցy��d�2C�������e���;���� �9E7�=sF�{�/g��h�?�V�V�����ʠH:O�$ꀹ�y�0�(��&g�Zar������`g@c�ry-#\�-�:��Hk0�9�<�A����bE�E�Y	����4p��� ���� ��o]J�gt�Moo/2I�X7R�7B"�������ɨ�y�k�*��J�p��%y�����j�Kǰ��9��7�u� I��=}"U̨R��z�>f�̕�^C�����*���nzj��.�)uUpȀL m�q��ݏ766�^�b���h��&�8�}b��dL2�7O��?��pk��D��^�,�8$b���J�r����]�Fn��ԋ�Fr�,���i���{}gڬ��N��'PO���};��{瞎� y���F�o�K�;h���;��B&����q��������܏���Q+��q&M��&qMVW�'4'�N���)�_L��]��	Q�x6�1��,�ϑ�9હ __���"")ɸ����E���稆%qy6��~�1�����+x*G:��KG�qy��J:��FZoq�c�Z��Tj�g�L+�bLCN=��T�9��isV�Cc�Jd0~J������}k�2�;���J�]�Y蕇%�� �P�Ŭ(g���v+�v������}��Q��P�ݢ߇��ֹ�Þ0K��	�E�[R���W͐�8����J���$Ob��j�\�1L�M8׀�k�=k.1���}T/x��Զ(W�j:��3�tt��	�A�L�L�V:S>�W����abҎ��`�'�`Z��U챞�����R��WE�_&�#����_�\a��[/X����_�O����h�'[�_�>Z|~�����
���ߙ9��Ȭ,9��5e����+��_�Ԫ=X�>�u��uQD�����'�楒=ܪ�
�|j�R�	ҍ��_;�Dsk(��ʎV,U4
��e'֐Du?Y��;���p�Mh�4�bU�סV�U-��@4�Q���˛�E��G��BG��D9j�z���~�c�f>�b*��I�0�	�+z��:Or@��з�z�H�������<ǧ���.=2�f�8���,��K	�ڋ�#8��?�yj�Q�Ry(àNB��J����q*�}$+*�k��%�?�L�y�w�|��.�E�@�R납.�/�JRx�]N�LKl� ��2P��=��t���:ğU*H���T>BF���__
=�Og���8�����T�q�&��iڼr�{x~����	~;�0%2���'l��V܆�5O�gHq>��G=�Fj��$�(J���U�v��A�A��s�L���n���)��1�JI@�b�X1�'n�z)j�Gr�T2����8U�@�y�y/Ո�Ę�������y��U{S�m����HW����/`�$�6מU�]��7�]��GH�_�ӡ8BH�9��FY�=�1g�T���w&~N��0���ۖ<������ >X�����r����09<e��i����]B~{�����]��_��u�u\�l����E4���� �[)}a�߳Hm+,R8�]�,��l����{P�o���N7��!�����Dd��o�:��
�*K����g�F��>��tR��x"�l���D{�ig0*��wy��aNd�W��Z��Pƭ<��e9lrj�$of:!���X�Ҋ3�w��.�L��Bv�4�x䗮�rF����	}�.xmMO�R�'���4��Q��"�h��?�P=���eYA��U��@���gj�7kc`���~�a֦N�U,���%!���i��Ew�\ڻ�X���p�;�,Y W�q,]�+���F6n�g�%*����߀�)�����O�����͂��oFÔ;ٻ�p���!L���@�=ԢY2F�?L��n������},Kl���b9�3����|ex����-��f	Y����8N�"�����.i�}�F��Z�8pr���S������"�X~�=6�.?9��lʑ��/q���P�U�<�����88a�s0�:bCιQIݪ���c�y�6V�h���,�<1��O��a�t9{��L�Z;�2c��s���M	�����R��IlZi=������Z�av���"����pn��,:EG׉"�#~rI��m��>� r���ӌ���A�]MH�qSr[��k3ʻ�u����i��DR�Ax���"c���XQ�z �ɶ�9糌@p9�����H/�0��Lݘ��A�XD�l���)@Pb��'t�9�>�7���|�x�µZ��,�T��=�Ai�u���t;*a�����m}%Z����yL���i1�1�H� �n�N���:�����
FTI��&Ţ�h+�NEx�nHC�|��0�:Go��o	�B��yr�Ո�R �|��{g��z11�;�J%e
�$rj�Iw���=+cj_:1�pVt�'�~�G�];�Cn
����{�v����C�PF�w�&�o�KK��@s��. �m�=�!_O�t`�ͥS��
"!_�º^7�d�����Tڶj�Q�%]�pQEH�X�3�L}�8��F�E�r�\b��Nͧ^@cO��mK�)!��W x/V������Ƅ��Y�GDC87Ҽ�f�n�c&1Wq'��{P7�����/�cX9=�����,�:�����һG�"/jx}�����&�2O�1�4�F�zJ�@���tY�����
�Ff��Ue-5u9>���&��33:fۭ�R_B(�X���A�+D������<M��L�ű���d���ǵq�%f��~�Ž5�>�	3{&�Gf\��>X���O�[����&��/]Ֆ�%~��/���<�gIM��|񙃁g�Rg0B麉>�n1@�>�������؋�̏d\�u�z�jx�nq4]��ҝ+߭Fř��-�9�8醀	�_��;��	h��÷;`'a�����d��pZ���t�JZp���2%��w�*�s���w���>#p�:�O%k�����-XM��q�b�nh0�h��z��{�r��k��#J�U�3zl
d0�C"��w��Ȏm����s�)u�&s�%Uzg���;�y� !��e��׷h��b�W�5 ;m�.2���K�Ͻ�d�t��#�Ќ0&�7~��>��9yZqu����)��7Ҩrc3�b���� |��v������1t���"8�=^�%��
Ѳ�Q*+7��;8܂s.��ИJV�(�	���iֲ��whn��醚�43�B�=G9KTƭ֍ӯ!�������q��߄*�����b�o0'���%�	<��E!lU�o�.�`����a��c�����҆�g���3��~'�)�͏��7���&ö��E&R���QIð��ux�����f�^�ح�����2M�����X*��юY-Pc�S�v�I����Qy&� ���ߖ@�k���k��A,��Z �F��#/�9�S���*��|q�-�"��y}�=�����b��Ȝ������U�����u�S��b!�,A��n-�����z_,Ic-�v���w�3� �r�܏2H��\����V~uF���A䟚�@�5e��U�q��g�z�B�ż��<�d2h� ?�����]A�ex�r,	|���o���� ��303�ڮL^G`��Wfa="e�x�0��	��X���C��j�I24�@. �y�s��9�׵�ZXn��
f�5�8i��쨾��+ F�S���~�5	[I�W/���9��$��LXIkBVPvҁE_\F���ۙ�b��>CNF�; �¹�P���װ��iu��E��4$���K�N�5��[
���^pI�ڄq#7�
Y��<O�{!�];<L�,@��ZH�s���9�]�Y��	<&��J�9.y�R�U-D�=��ɡ�$l�j_�f�H�e�UQy��D-��izY�pk�J_NX~Z�+�(�B��!�?HE�M�>��ż>K�:�L�U*r2׬4<f��{���]�`C=��~�+�F�/.Fp��tX���Mh9+u��QM��P0	����ʵ�x��2��L6��"T�U论DC�ϙ�4�p�ߓH�I�^6�Ï�3�����Y_���h4�L�.*qC��;�����)�0)�s)F�$��l��
��b���sݪ�_��S#�"o<�$>��ٹN���I8�s�_�2JE��{�0H�D�^�[���@��$�-�P�g�1ԖV�\(�0��ͻ��i��0�����s�y��|*�)z���籔V+�E�=a� 7�˜A�t���;��%�c,8֔��n8�i V+x?/dp�����J�/%���z�Ŭ507x��H�r�{�<�M��';�v�6�u����6Q�
�����ߔ��Zq�Ƹ�o��wS`����#�&4��#��1��+E�w���1dŎ~*������_:�����&�Q�#��C���:�8�N�Z�#��1�?��J�6[w�<���>I���%>��=5N��]3H:'펿h�N9��+�3�-"�,xm�^ᾎN�y��|�W�;�J��P-�!�kV�2Hi��Vr��p�*����&�߼j珦oB���Z��T�OoH�{զ��-��(6Z9����v��bg)��|ԯ)$)�7W�u����H6���o\d��u��7���*�HZ�30@~�������K{c���}ǹ�3�J���MX+C�A���1Х��dT̾�d�1��ϨQ
�>���+�˼�3�I�S�
9���瀴H�f:�f@�D|`du^���uX����lh�5<3Г��Q���%�q2K�g�<��"�=i�7$Qn��A�Gך��N@X��
�g���7˼eҤ�m���N�g҅��9'��E�_7Ĩ�D��W��睾T!�{�8~؅33Jz���
�|�|�i��3�ET�ѝ�f��G�}b�-��Z���&.��{��%�wuv��?*����_]�,�B�Om#+s"�����̖1#�� A�N�Z��TQ��[��l�[�σ)^SKg�K�f� 0zBm��$��D]�O8�( �;;��yZ6�p*�i����h%k�r�s}��5�`T�"����*�I���E/P��q�\�bEN	?�[ԟ����r�Y!]�;�i�)v�+v�_6]�L��Z�=:'W8��y6�!���y��)b9�F�DWҳ����`�h= ��GݷS���o)1��` 9�8��F�<��nM�����?�'�R=�c�>�A�1��2��&p��i����!���z~�P\,|=!��InH�[�����Rb�c"��K��v�<��NH쓻%����5��rYy�6�n���uߠ��a&<N��2}�s��d�����%!��aW�/=�cg���;��]~����>��h�����KFz�����(p�8*��!�P�3dx�c�������U�i�E���p�ͱ��U��ex�(�i^���׋��eO��{Տ����ci�%ۏ:�5f3AP��oB��b�Y�	�ڷҥ���4��_,Buv��ˤ]���Z��$�|����$��;i�����fRJ #{�����߷{������u�`��E ,mR�Q�� ������������5�-?-������S)��	�i�;�c�$@o�O\� >��Ȓݞp�:~Z�������｟�\���$��o�������M�
��%��C�l�",���F!�r�N]K��D�i/�-P
���]-K���#��I�cNi�Esۚ@Q���[����H��eZ�cݝE��qA�8{MA��{��~.��`GgLv�u��/M,dx�5Sm�
y������q�K (�j��.-�
����_��sZ��1�30�X��z�8ߌd�q/���+s^07�i<��gy�bm��V#JA�w����ȿ�W���M�m?�
��«Qӊm��j$`�D&��cV�i��s�[�1t�/�8&����b��Ϭ�}�:Z�3���oi�]�D�Lv�(ɠ��������Fvc��"i�!FM���O�>5V�f۳pi��/�݋��������rs���r�6�.��&�9�G'�����9M��W���p��$���w5W1���
��4�rR&d{�;�D#�B��$@]vH"�6�V��ڬ_�-`�f�1������Zh��EbU\<��f��":�.j�Ql��J�m?���N���,�7�\�c��O������Ͷ�wj�lp^��$?v�G�@���(�6�~�������|XP<���Cdr���������V.ixF\���~�-�,د�o�;��=�l��C*� ,;��+����H'$ã1��`g�	]����d�|P�[�R��+��n�6���BZx��^Xؒ��<l�]�a�CV�\���(]���*�Q@g�T��w�S���#}�� �_�W���o-6�q�9�t�`����c�L����h�/%��Օ}>����`�#�[���Q`}g:��,�m�[	���[����`1�'�.^�j�Y&M�Ix�=�-Nr�IfQtM�᤾���2Rq��U�6�����؛8|���|����Z儱���pՠK1�Mh�X{��0	ŉ:�ٵ�e�/v �ɭ��p/����΂��$���ٞ1��;�պ�p���ћR�IO�θS�?�R>C��O�C0���0{����+P�H`|Q�O�����&G��r,OS�?4�4�vbݧ��$�Y9���g�|d�m:�ٖp���.=�x(�Z~OWhM-H����s�"2/��� �L��w���"=�r�.)���T�0�g����
k���<Z�����QmF�G���f"ɀ�����7��i�]���ۛ��j�v��E`�P�Dq��Ub��"�+�T�Xʮ�$�7R^JEg�j/@侗;�!�$��{�R����W���D�HW��Q��5��&i|�$��uZ@�_��h���'Z���	,�p��g:ckj����<c>������)S�6�m�
_Zi�(�[��}l�@������F��W�{%E��Y{0N�#:g4��JY�t����^&��@��I�i�h1 �bd�6�I� ��IY�1p"�Jt��Ք66Vj�7�Bs�	��*젶&���|��n ɤB�E�^IerEr��ua2�e?���VNP1�6�n�#���)P=L^tD~�sTmG�����{"���>��M��Vj�邷��,B�7T��'��8y�)bs��1�yS�J��6�;��+��6y�{/iY3��-_w��0D����^�T T�
���sV`��k*9?� ?��]�F����B����*G� �*��}H���Nt)+�W�����R�~j,>Kȏ�X���h�����
ܝ+4�(��R���{$'C�%���eQ�BOӨ+(�}�k����*��Uc�n�a��|��~υlRSM�v�G<^�U�(�s�_�B�����XI��p�|�U{�)7&&�O��+ާ�{�[y�4�6��A�뮧�h���E��BB�^�RF� pK�g�kP�N[�Ys,y�ds_��|S���^��|&^�����^�C��C�E�Q�ǧ�d}��_e/v�h��nv��p��8���5^x6�Wzӵ��^�^"M�$�O#yc"����O�>P��[xJ$!�@�q�,	����S�'П5}�*��1wݛ�Th�:L1�!1V�P�I�����oW���L��{rݰ�����mE����Ix�n����+-a'���t���k���P\Em�wgor�����-ÐU}����
��1gȄ���P:��H�RT��m��O_�~���k��=Q�2�
i�쒛��=�A�E�t��)���Zx�?K���~-4������;��'<S�S�L�}��9���[kJ>:��N�����(�\���x������7�c%;�Jֶ��O�.�vk��(���"�`w���y%QR�Q�Z^�=R��2��c
���K��	b��.��wd�lR/?ъN�T9���t���W���'+�|�^`�U/P_z>=���=Q�ʵ��:/�������p���_�J;z\y�yC��jO#��u�%����'2*_C5�6�g�%����U[����+�>(��*�^��CeZ� Ze��҄����Ư$��j��r��;�:�[��pRޣ�M:pĀ��Z<ofd�is/�k"�a-{i����$���|e�[c���>n�����2~�y�e6ewY<wV��OxN���:?fR.dؼ�JIi�O����QջӪ���E�9{H��y���~���q3��, ��X7Eg�+���0$����=�� Qvܧ-�I������y��:��#�k�����ރV��FQ8�DB��g�oPi'�I�]y�eJp#!0?��B.�Ϻ��j�{ĉ[0��I��2N�z����(*wWҧ��d;u6"��f�������C}=�̛*�1�_v�w+#%�$��|:᱃����
�FUvT�"�O16L�N��r
����-�Ԫ�%�ő�/�ܞg���k:u��j�ç�ȠJ�r�/@o2_�n�$̧�_�*��@�r��cEv�{�<K���� �'�aN
1b&H~ļ`��"=2���o����`�$"L�X�E�&�vD�O��V��ўq2��x�X� �JEμ�0oUo�7[\T�Y��tE%E����5�1��n��=���"�mC�\�͓>����lE�Cd��]�7]��hwK-�!�V��~�Y
3p#��v;�����v����"��ۂj���K�e����6V��{sD�Wl�t��9�F�����6�ciJ�ʖصBV���qJ�P�I��|���6���SS��]X��i�J:�0\�LrB�x�/4��ɡ�?��ma��[<�5e�0��C|�`㎳�]ZA_�;��GR�d� G��b���(��
��%`���T�!�"��v!b���C%F��v-�|%��49��'\�߅��5�������[�x�p�Rs��!S�������B���kY������\�}}��&,:�s��)��1�*��*SB�O����'Oy@S�7�p�I=)���F�C��~2J��{Ӏ��(o}{�3E��d�N��D��{�Nf�����rt�3�����*�n�L����+�$欓���a�F��4�� �ČU0w�&�Z������=���sH!f�c��.�]�7��!�����ə�0|������۵}ꘌ�����Əߌ|���j�ϰ9��-��}��Z�+
87�X��C�1������������;�q����J��cQB$�JEDp���z��.������~�ze��_ڀji��3}��{��R�&���#��	����o��݄
�Ue���f7�}��5>�t:����]��"�,���<o��q��J��vw(�yB������J�%a��+��*�@��ſbgN�]b6�cI��2��"\�j�k�H�`����B`���?�O��� hrs��2����Pnݹ<�b�Uӫk��0�]cs�f"//�[=FE�j�л����K$�L�yJa�o� h~M��F���j���u�}�����\�ڮ���ų���]��/p��r%�C����x��0O����^����J�� �w�0�]%6������9�}�S!5�  ��p��7YR
&}ϒ�É'��>��K��j�Ѧ��=3��G��uu
�CZީ����l��!�ގm>��ynВ.�ƚL�v���
kL��?�+���6S�`/T����{ 
����V�1i�.!��b�}���y��<�\�
�&�l�)�-�߯��Um�$)�"v�KrrZ��b.�[Ӹ`[k3�α��C9g�	`K�r�ׄ��Ր��"����g����~߻�s>8)����9���Aao�Q;T\}�UcN�黏2��$U/	���/\�r��%�AN3�/g���u8�!���m��Z����>�r�.�O�l��46�[�dB��������z�	�Hi�_�숃k�`��D��^i�
_rf���>B뾴#�BZ�?�鸾����Rbpg���f5��݊�w:��6{�"*b��Y��t��F9W����W��T�|3"��,���dòY@<�Ԣ
��0a>�k�4�N¿2��@c�+�LU3��� ����I�ԩ@�?��G�hc�;ᘩ�@QϬ�ݺ��Q���e�I%6ݓc:MJ���[��_ik���5k�J����O}�䧥6	J��Y�����NB�w,�^n��)��mP�g:Zs���N̄��[ue; ��5�X�����O	y�b�<�^{8��~��}N�-��l�sȆ%���c�q��R�#���#��fAw5�l5��T��5-F����J�������`�(-�ZU?�6p_���M���}��Eչ*�V��yB��S�s�wyK� ��=�nG�S�o'�+	K=�n���k��� �u��=��K_����Oڦ�WS����NC�Mwa���&���`!��4�W�;Ry�f
C�-��ڗU�7��B1�xS�V�:8)C1
Zv9����&�:�R�Cp�`��ÎC�)�Y�4q����	�{;0�1���qRwTP��E1w׫� u�����O�C�G0
瀆��j���bOGVB���M:-���}��fߋ� �.��^B�&F�t9mF/y7��y@c;���E��ll'8�b�m����x(bJ�|(HX��9qٶ�;Sd�����
��F�C�+wx�j`o��/ڛt��X�
�B{$��l��TB��q4Z��JsWۺ%�����Q�!����Yo�.\�4�I��8lO�~�Xi!����Ӣs�R��L-�L$˺�})E��N��1�%�	���6cK�Cπ��&��&�,?��GB����k����Qse��5<]�`8��=�X�%i�s�򇪐�}�H2u1&�7L瀉gv�X*�-T�\����`��̗G��Di"v_o� �v�~�'��߬)!;vKs�$ef� c�#%Ox��}P�B�Z��4��(����֚��O.�u6�e(��I�$��}�$z� Cܔ"��P��w�ёlN��6y)���`����:Ff�Q���k��������5���)���ɍ\��Lv'iz/�1 l��v��W�wB�RQ]��(�����CcAͦ��\�ՙ�K�/L�T��e}t�ܖ��mLQu �f���Ӻ�9��g	�ep��](T}�-�K��sX�4�v�ĝ[ �0��=��)A4������+�E=��	����q��;%���R�aɥ����fxDX���ɳlmP���;*�-�8B"1δl�*�P_�6�ld������̮a%;A�z�Gn���E4�%r�kW��H�Jg�3K���D�)��}�ˑ�Cӎ�����Q��)��Sݎ3���^�aLْك�5v�d��%͸�t�Oټ�"ï¢� ��~�|�p�Z�<
��ӤJUa��5�p�SJť��f(˗�o�ar3�M�.�j�z��0O���D��R7o�ꄒ2Yt��e�mkͺo.�%k��n���k/f?���Y��>b�іMa/����oe���Y��k���6�R��)�R�6���Q�-��t�h}P8�u�x�*�,��Ó���%,��������v���A>�vK̙����.�zmW��>����O�1�$��xHG Vu7���d��)YI:���`)������u�#�-��$B}lZ������h8��q��f���o(s������Q�6&�{�o���2��n ���qW�5$���>sOM)Aɺ�a�}�`�s o?X���|��h8�����8�_}Rk}'���h�~M,�9�����-�L�YH��� �"a�\���Q��M�|�w.��A�'��e��5Î��$Z��ʖ&�w7�'��6K���@��\��N�n�؁]'I���Q?D�����|p`����]���[i�:Q�f�����w�:OC�%񦬬!<���Ā� �@���_���Q�H���)Њ�\��=s��Vj����)?�Y�Iވ� �c�+B�wq���Tٍ���FS�$�n��C^?b�}�y�>�INvz���?�짙���uT"�j�J��!�c�8'�K��h�������4/i#� �z�"�o��4P��|��[�x��������b,2~$�[h�_��r��!Б ����An;	���kU�a���<-��5�G�\l����R��I�B�j�v��7�T�FQ��o�A�D)q����nư��Ut��_a2Y	u=�i$�;����)"m؎��F�A���K����E}D��!��w��]6���6����8y�h����h���^ ���l�Ѳ��W^F���� �u� ��Pb't�b�z�)��>�2L-�`k3g��.a
F����e�鎌3<,�=,w=Z��d��U��.��|���B
�ֿs��l�@b#`��~�>\���Fx᭶�5�����?�H��6����h*�V��~�\E��}�i��"��Y�x��:1�*������`�b���V�h��$)>�`#43�1�����H8�5K���~PT}��Ԑ���Rm�.���5C�LhW`,�>lC�t(|so�2VU+��Nע�b��+"6�Y�p7{��G��L������ذ{���S��#Ȝ��?D�I
��T�����唤��י�J#3R� ��%p��,Nl9�*��Y�])�k�V޳V�|�����tW�T����p[�XѾw���M�Q&��^�Z���0�`���QNGW'��DM.>��Q�TSO���V��U��(7����U-���
1(����e-���ll^k��Bj]���j��/6�km�H���m���40�⟃:w2سTk�������������4>��䘏ǒN�X�nT �i��Q����mCk���F�6��qOn��.��'/t3�6���	��c���F0o\��[
����e����D�R�V�^�3��>�N2����pD��\�6�aY  DO̡�E�6
�nqLDC�Z8ɍ֊T�?=���57��{�\1!���������(��KJ{�YÑvq�2�Ɲ�4�����H窆�,tw(FH�P���Ѭ�R?�r{"�j�{ �>�scgKi�4-�J��4�[@5��O�l�U~��|`#=Φ�o|�����5����综���M95�@�U���|�,��|�h����@]��[^n�94h�E�����KO��F���}�\��W�cf�=��_@N(��D�}Z=�g"��L���l'�]�H��砍����l�(�@V���EA���J_����W���i|��H�(�d!���$�G ֦
x=	N��Rqw~ڰ?#=s����K4/S���}�PFL��W���PK�%�]�5����y� ��S=چ�%A�1�u߽�V|��>�NL�ϐϺ44�~x��wk�^81_nmU��*0���\�l�ovn��n�t��p�ҏ
�dį��ݵ>�����f��UA�����6FN��n�N��<���V�L������37�p)6NF����HA"���"a�/�8�Z�X�F�	2p/5�\$�\�c�G�F��H@�[Hß�x��ڑ�(8�1��L��5�P��QGsvB{�jH݈�S������FÜ22% `��9`�aJ�{�뵈���h/G�?x���T��R��D�@p�a*�*��+q��Li0T�34�����]��j��y�Hw�y��4LMӚ�M+�R������-�:A��I��@G%pH�aJ�<ˀM@�	��"�p�nt����@�vΐ�fW!Řm�~��v������ʫdH�����g��|W �9�O�
8_2���݄͢A����{�!o	x�䲛&n�,�ot�����O]�y
�UJJ9�ڈ�}���eX��������G[��m^��y ���_"����ZEY,X�}���El��)�0�w&3�[����\�{H][�9��g����w2>05𪸨��w���ttO#���h@�}�|җ�󎑍:�"�K1j�q]�����ε���F�	���|}���e�a���������dװ�Y���iB;�Dʚ�ՑGLx
zmQ�Tؼa�u>d���;�8c������+��c�f�A�!ܭ�*�1�qc��W��{��O�*g�d*o����~"�,�$�v]D����
�7н����/^�y_�".�K�F*B�����z���nQN ��ZH-��A3��i�jӋ��.B#7�4`�Ʈw�\E�[���S�Ŏ 柤������zs67�H�ߜ<2�H�8����E�R�bº5�V�^m�i6ԟ�rۛ�� �c8���n�[;�Zr�����
�Y���G:��>S��q�� 9ϓ���#;����a��C-4+�̆�x��(�����q�ğ�7j�t�=w�� k���tA��Iw�RU�I�P�h��bz��S�n���i�d�ڢy��ޑ�	2���	�p���Զ��-���TR�m�I�=���R!�}Ē�<��%�Ey���hZ��`�Tn2�>į�X߳#]�O˶����ȋZ�0!�������J�;CB�x ��6�v���υ����s���S��츇���x�+۩ݲ��x-�$�O� #��"q�>]R�n����:�9w�]��#��P\J]���(��I�� CAW��|��g6���jK�G�h�|��d	)��{b�i��Ʉ��J^��2���ՔZ�M�(l̯0�*���V���]�{�}-�u��w��S��֭� �!f�m���t�C���e^����[���2��S�$�
N��Hc�%��6Vq[��C�i� i�U��:����1m}d�fH�f�l����V0<�"8`�z��M~�vx���1{�ʮ�0O�C����-�/���:�3k�D���	�n`��C�ԫ������#�D���~�ZL�b�q�e���3��b)�V]p`�YM�|�kA����e޺��c�z僼}�G��;�}N�3c�%ĔhS��vNN%5=�L�e�
�09��{���&S�xBUkW쬮����;�	z�J�׊4ך�.Cv��}���LfdT�$���k�q !?�b�3�q�j'��=E���D��]t�3���ۦy~�<;��j���Ɓ�*7̡��c���0���0���0q*;�nב�il�D��N�(�/�o���V�}j���ɿ��Y�(���|�W�{$tГH�H[FC�i(����ʒ��+���+C��
z��Ō�*l�un����]��S���V�1%(�ZW\��
2~_��_0T9%Pк�"V�1؍���H �*[^�7x�*�����E
��d�������̚6��ˋ�n��
�<�$����%<g���2�x����"��H�ᨌ/Թc�b��>�j1���y�z!����vqM�-�l>��$V��PS���	�P�4�:F$M�Uz�˜���eK7��'.��N��@��X�S����-�q����߀w��h)PƐdi�]��_���"�0nyC�H �.e��n �v����u�U1Qv�86fV�X'�i�.�SL�,p�8�@;��<�L�&r��w��)d>��ӓG��a���(���2��a����=�X�<|ߞ�}����y�~um��jwH"�X�Iץ~�K�BP���$���`�v��?� S~��l�������Y��/E�F�
�b�>�
B�6��/˷�� ʊe�p�����{��D����ٽ��:2��4��s/ ��o��c(���b[���Yj.]���b.SN�k�?��[n�����sP0l�	�~@H�B��+pm�WhY � �w9��(j���?����9��/��h���'����-m����S5{���J����ʡȥ=��ސY�LK�Gz����*t�nF���N���Rx^�=�5c+?W���J���>g�h��ST֮��1J��V��[�e�V��O��$����{��/��x�%ܹ��.1f�Jh�P��_��w%�5�QuC��:��b�6���@� �J�4��6>��~�˴[�/�J���&������Z�?�ʸ����DL8�5�,��|�S}�"�Vu���Ϙ39H�eYA0�~Q;WHK� .];Mf>b�Nu��7�:- ����q�����UWK�ѷ�Z5X�;s��xף�~u��٥�U���9_m�ZK�#�?4z���%【5 �q $(?����Aӌ���sc��f*1�d�p�];��Fw�����9�Ǳ��iz3"غ�HNe��������g7��ú�#�x����/���fTh�˯_�蹺�s-����1��3��.+���Q��P+���8��x8f��7�a��8��,�`�a�;�u���hl�^V,��{Vѯ@�WJ���L`�d[t�9=�Q�c�Ll�=Ļ6#�u���Q�X��ae�O�H���F� �RI���o?kx��#	@�Zz�GG�2;J5��%��K}�2�(����tv��}D,�঻h�}h8g��_;M��a_@δ�~շweн-|1�!	�=lvd�%�%h��n)�of��#4
~.�y�(�������n�m�2������4�MGf�V�KID�1�!|ʣ#��J9X�>�CG%
[�]_l�,b���;6f:�h�ߩ���[3s�՞��W�w^E���z����jˈ���5�.Z���'�2
V�y�o}�d����*B`��#T���0Z�j�!�U�>m��s�"�t`p]K�t����3\C��<��٢|H܈�	(��u{����8O���3wɦ�=�!�aq�Z݄�7�ǫ�x'�a����8��<*�]̶� zx��Y3|�yi����Q�aQ�P������*z� >��UY�iq	Y��e�� M����wRX���*�8oy� Ґo�F�F�,,1�`��Z���� ,T�y����n��<�3e�SA�Cnu`���q�Uq�9�0$vʴ!�m�8	Z�Iq����t<�5��BH�QY�!<;�ٱ�����(�S�%M��GQl��P�v�9��U�t�f⒓L��hOd���9�G�ֈ	<�r��1R��r�-�i�堷up?���W`9���I��a�nM�0=*��!Es|hӑ�n�c��!��ޑ��X��f�-sWq<�������?����)�������'gݎ[58�9̯-1�gp�(�����HP�K��\vw>R�@�8;C�`dr�%7JR[M��9�{\��z���r�`�	��w�n��秜F8��i�mZ�������)z���gi��ryr4%��|!�ʱ�kK)#�W�B�T[��P�*ל��c5���Ww���|�_{�v¶��O��g�x�$_X9YSj������F�QSԿ/c���A��Ψ*A���@����c_�fKB��5F�S�p
h���5ؓ)Y@7�ع���_��d�Bav�{���fD"Q�_o��`��n�N>R3��y�����/�c�5=�(��\�����I?(䮪 j�Uѝ��U3u�:��-�}��ӷ���ܐyz����kV7���	n�w}7AB�tY(aO>A5�C�؛�1�_٢Lu��I�Otr�P��l�&�&�7��i���Q�5��㞎��(*�$�#h��CȝX[=�8W=�.wۦ:�{�{/��k�k�Y��3�9�]\!�U9�O�3ńu�}�(/`�$���0�e����A����ruC��4���٣F�c"E`��	ݘM7>�Sr���B֐�\����C�R�L�֪���*��`j�/�PKR.2DV6��s�t��s,�~��y�-��#;ό0�Xٶ2T�W�����0�ȝ���@�ph<�f��k 톶s��A/�V��$�8/=��Rm�-�a8���^	㿪�>�9���XM>>�\�������CӭX6��+�N�,q��wZI�u�>��\=jh�-I߈������n�2T�ØŔ�&���]~ऐ�.a��
h����A)/��">���9A�/0�,��]H��[ ��(�ch����<C�;&�zI;G��;Rns�ȩ����	F��ZU�|AyR5�P���ړ#��;\J3y�<�%�xB�J_�4����(�,��TR|ػBF����,	�˟G�FlV����c��Vt�{ik���S���r)!��+Ђ
��D�����g�M�[#���fI<���ʚs,��#��$�RD�?�÷��ߩO�B1� $����#7�B�n]���`�ʆ�����G��V��g��~2Y�:@T���ݞ���ٶʌ�%��D:0`��u�f��U�7��mƈ`����|p\gQpy��ћYU�k�i�����=������lEXs�KcVw,�.0{�k>����ɵ��)N�q.���f��F���X��+����hWG��BmK���z�̍m�0/znS_�4#yX�\-���u�y4Ҿh�.�%F�>���J;�!GG -{\�6�&�V�t���i%�d|�}��gـ���Z��D�����L�<�KN�Rd;�z�xV#i�Vt�����_��u�픪��b��%���92l�ov^�r�4�1v�!�8M�$�+�7�.�����Y���~�Xͼ.�E��5�C�@�ڣ8���"u��'J}�����T��\�	\�P��T�N�s����BJ��,�:1|MV��B�Q��{�I=U���yB�vWOFKDG-��N s�]P��
���1R��9
�����D�\�K�����oŖE0m ����71���	|O���LZ�D�����VZ��0�\[�u�Ϝj�}���7�~��a��>���>���![�(����d=Z�q�p;���&�]�7ܲ����\�x����EE���yu/Dd9~K�����|� �2U�?�P��n��J~�ȕD��{����0�w���P�9�B�U���	��
�6q4��w�S�V6w�V����r��h
�"�/��mS4�i糞�d�N��e�K�V$ �lo�K(�����T��H�d�����&2Pz���[f����UR��x1�\6��q\f�X.�>��{��B�A'Q���0oGX��D��{=ly���&u_����Ζ�HN%�o����u1۾>sg�ȋ3���HxA �i�ײ�ɝm�F�I�ڧ�fx���1|�a�y�ܜ�|��Ά�V��xU:�Lg���ч��x%ј1�%WY��=�LK)�X�ϙ��c�Q_�W�HA�zat�ג���`��\4m����2a�y��a���_*���ZB����	����'j:�$��v�n��J���H?�,6�p�Z���F��)yW�����!�fO�Q�<3t�hz�W� ���Y�L�8���.��>]Q���/����;"�w��n�zL��|�7�Eq�W˨ �}�W���p����ML�"&;-^�WK��H0�v�K@�U��0Jj�8�؟q?fmm�|��}.a��@,�~��a�i`�5`r�4Qu^��k�#f���Ǉ����Б�=Jl��E@R�#'UMd�Ag�r�-�Qle�o]���۟����>=��k�YT.�t�����EIni��!O���g�MWj;���gs/"��;0O���\M�Y$�� Ս�C9�|�ap&��O)p(�'U~���� �I��	�r	����h�s�y�}���w��c���=T���Y�w���d+u%��[	�����!���g�[��\�h7����c�I8����ur!���)�����퉧a�~<r���8�O�dB��u�%[�3Q�L8�~�dye��_�	v3��T���f�h�#L�+�$��8x3�B���T�L�>��u�P~b���>zG�n����n�a͗h#uz��x9r@4M �j��`�'x8�y=�-	�!	fa<���1�]L��g�qv�⬁9�X�c!m�|f�??~ǟ�db�	�"���[��K��i���M���[+��ʕ�i%����g��Wv�6����њdJY�n����p�T8ϼ�T�̆�ƴ�av&�Z��X����>��	�82Y��ŉg�\��H��J�`�P�r���7X;%���x8�axD�ۭ<5��8��H�+���O�
v֐)����p?�./�OkE�Ty(�𾨒���@������\�p���q���iMsr�Nr����72��5�Ǝ�a񏛺0�V����[�S�e�l2b[���y���><��]A�hd�P�C��DI�b�s>_4�v�J��٠�΀_�5ri����_3O���d���Mv��Qč���?R���L�D���������fi�pě�J9I�J�M�b�b$?Y�pT�����f����.�Së�*=���$��{�����<n�>�O�9qR��.9�k�>�=�d�t�k��MD���_^4
A��k���j��}�y�J7VI$����Y��ɽ���ֶ�+B�:4%���߼k�Єl��*<��O[<��:�b��iCvB�bb�s���@�H�Z?˸��kQ� ��m}��	*��DP?����Pf�5R,�"Ij�x�r��$#��~���S�����.Wf�k��Huݥ$�z�.�&�>�J�V��O2�]��QO)3�Dw�����2�it���~�7���^�*d�=�Fy�֘f������1�����}�~#Pȇt2^{��f1(�F
��}�pN��;�����!6�$�V�CX��R���;H��f9��?���@/H�@,RԆ��q�T9�� f�l���U4���l�dj%�ϛ�7�Hݯ&��'�9��_� >���i�]�.E1���H:-��n/�`�E���
��߿m��]��P� u����%e�:=�ڨmB�t�!�����OXs�Gt|u�������6�@u�~�O���*}��}�[�A�*���i�5VÍӤ�D���C��+�Ō���j�����<�B�AG��՗��jS?$ph�10$e�R]:������hZ�B�pA���h@�XL�Q�;�jQz�ݪ��H���533���k)�]x�/�L1�͓ŧ*����ڲY��h�.�+=l��^#+���i	�R�
�^��([�Sv�Uf����y �<לs�.�*�۸��lX��/L�o��<1({���"����^~��Q����h�O�%�Ո��Գ<�~�*��1[�{m9o��y��a����o��#�*~���`*8�s��ݐ��a����5��0[Ii��:N�H����l��Ī��*^�F��e]�{mh��!��c�*l�I��v��jѮ����4	�RZ�`�����,�z� L	O�u�}�h�o!}*;���Z|Q�]�[{��g4a�����]9Vr�6��A�#�́���8�S,��Hư�axN=�hLSK�v��ݯ��M������٫�	M�6+&��)ɦ�2D(�ѻn!��с����K3�%'����m�ú����&h��O	��������~U�#
�e=-v%�=����>a��`�0�i	[m[l��1�d_s�0�8NӁ[�R1jz$��Sa4v�q/q���I腛���+DiI�nr������W/2Ge�%��f��x��9Ƌ��
��8����[����j�"�O��'^��j~�����`[&��!M�l��$��}d�<�$�V9����^�w��Gc3�\w���(?��DK���'�r$2��n!	-C[j�Y��:�t�f[x$0�xӤd\,�m�n�k|S$R��Ρ*��������� 3���5�.\C{���l,��z8�g0kڿD�����j�8��Ts�Jl|]~�Nfʔ^�hK�7�\�'1^W3��������nh&y�7��z><>z��p��j*8T8�c�d�zWR`߰+�7G��c�(7������D� �B�$Vke���Y������&�:�}��.��7gQ�sz����Яh�~.��q	E��%��g��-�����V� K���s�Mkf}k��/�l�EE�{V�t���k���{9�/�����#΂�;{���f�}�C'�fA,�6��_��M�!s~�L��bי�*��ߩ�c&�1yn���N�oK�䎔9҂O�W������S���ˏ��7�`�))���@ʻ�_�I;�V�2r?�ĵ���������HS��HVb*��$���� �^���+���L��2�g�-���[��U�}YI���&wgL�ΙwŔ%I7��x��"Nk�A�'N�O�-!� ��}��M�cW���>S>-�=��P"�A�Rk��9�<��Odb8�(��/1����z;��V�I�`N�����f�س�)�k8krt�ZoGi@و���𖺂�H1[s!7��8�e��QCM��HK�W�4I?��5(��}䕄��D�y�ݕ:�	���0�g����`C �(�\j�:S̜�ƽ!x��^nn����-m
��I�Y����j���D+p�W�_�����Qo��/L�	��cZ�'�%ޔ�m�����w�j��s]���b�-��"\��A��Y�^����טyE.� 'ڭ�]Ǯ��8V�_�v��G`iSI�zkn)�v9�񏮵 ��U������=�$�$s1 �z_-�����e�d'ʷ��Uɖ��Q�;U��b�<�@�=Lo$K�� [%����˞���OH	�jU����\�����8��<,4����C��ki�Hc��PTz����$����hq�s�u~Lu�H�ۈ����&��T��� ȶA0�����;�\
tÓ�~�-��Y�~�h�7:l����B�i*�c�QL
# ���s�gU��M�����ZW��&u6�fce�4xV�"%ϲ�+�	O�N$q7fu��Q�"�1����Υd^�|���,�NXn��E�l�C%��ܡxΣ�9�ɭYf��;n�۩��Zt����l�/9��y\��fnk����n1hy�=G�& F�VB���}�%��f ��P��
dXO"�����#����&�����ߍ���dXÒH�� �O�5��0�S&�&��/e���m5�@�>�oP�f!8��L��ż��v�tj3�2޻	8�r�
��U��f��g�#��Y��/�ʽ�H-�9ۅ�	��N�*[��H]��*���I�&��<��4�َ���eW��R�����{d�,eWcDe�䯴 D�&��w� ��C�9m�',Q-���I�s�WT�?nwn��k毷As�̉���#��v&�^��{.i����y!%�{���ۏ����@�(}��Cl<�~մ� �B�+���)]\��(0n'_fi�e;��B+Lr�y��(&�MUو����E���?B"uG�;C"j���L@��섘���pL:ɆԆ��"��{�֨Υ��}�(`��+���������T����e�pd�zZ����{<\yf�%!ͦSS��k1�Q%���B�kC����!+~�{��;ow��|�ƾ����e$�`����֦i�la[6���_��ϒ���D�TN-a�N-q8,��<��A>����̶�P~ TwZ��䌆^����X@��n���7��޼F��9�j��G���ẅUiGfN�����:��	����7�H��k��89|ϰ|���'X�l��KR��2��G�^$��:y����ʾS�5DC�`�BQ)Vݠt��-�sV�D�
�,�B55N@���؟G�� $�8� �X��Cn#��V#�>"r��c'"H!T�	�rл������q�J�w?�²i+X*N�#ѩ�1�J۶�d��WO*�Nz����}��ͅ!˧�4x/���[/�k{�'���4�x��k~��9��I$ Ø���+�_M`�6[Q�=�R�O�%�3.K�5�Xh���}�[ꓩ0�+�I��J��S�%���[���/�Ջ�Y[4�w�`�s�k�5�
�������R=Y��C-ѽ��b�'\ ��弦�A5�⠨	�K B �����%t�y�w���������gѬN:
���^�Ώ�ߑ������a ��L�/0
�5����]#5u�#^v-C��/�|f���b��R�ܳ]��*7f��6����i�x ;��`��䳬u�,
�;�oBA[��S��e/��T�i��\i/��l����[�Q���%p���+_�t_T}����i��~�M9~ծ�ʶ�C�L��M	2)2a	/�?-V��|��<������*���i!�W9f7x�CbII��׽����)d?�g�QWU�a��1��ܩ�u/��B>�{a�Kr��+��O��L`ڌq��B%\bD-W�f�^�LDP��~���Sxd�buM5x�9is�íB��>�t!r��=<-f�;��S�#	���8�����qc`�g5ur�E��_�$�^"��Y�5�(�^P�H&�-��r���)�-�9��-+{�t�W�_;L}\��I�p]���}T�O��5ةD`7�8R���U��J��"\Ȗ9�=[M'b�g�U��h��2����n��E�@Fo�6f�R�ޭ�@��7���_�]顜%�J�g�<�67��w�ͅA�4��"�z��vT5w�*f��*y�j��al�i$<pi�s��	�"���3�am�Y<K*��]<��C�^��.v�^����),(�b��t�[���լ$�K)5�%)��伕�[� �ڀ�|�E��# �E7�6�솭�����1dRQIUx�2�.0m��)���pW6�Gc�}J�ׄ�(�T�'H��;}"VU]�xY�4�:�Q�Ȥ�Ȁ�@��_�NWS���h�.����f�i;�1:o����E1+�b�^�jc�WX����'�ءxn>f%n�D
�t��O���a��T~V�-�=��������l\g���VX|��0��f:�45��5Svu v}�J�V�����rFwͶ	��i"�0���~/N,�u�sl���ɮ��N�+�ں��>ҽG>l��i2�@�z/>��C�\�z��SR�_�.��1�<Mu\r��IW��_'���cS��u��oEy���9$������Ӓ����O� l�@�#���`��t��B�<W�o�&*|�Sl�EC��}<S�X���͜{b{��8ai� �00�i.q���˻�
��ih3���4�j�`q�� `coI�z��߷�X���������%g{�Emm� �J�R�H���l�~�D�V|�Ҁ��KH0�T���s�2�]�`��@N%y�q�=�܋)C�|"��ř�҉�A���Lđ�� N�����KS]GX�� ܵZ��mѲ+L�۟\l�-@9 ��Z{b5C������i'%	��	r�& ���5�0��|}�2Y9Mې&�h��T�u�%[܂�s�A���أ�W�,�YN�'�k���[�`��P�G֗�Y3�BB�����tbH	�1�1#��
�|	��/$��})eGO
�����	��q��ɫ�g��t#�Y�C�]��7�f���N�ޅŖư��*��؜��-������*%���/��č���)lS��B,�=���`��E�d ξ��MY+![uiZc5����,�N*�"��=�0C���c���ip�C��{�͖2���SI�E\ʊ��� �W� GՖ.QQ�枖�oi�~��yE��,k	���1f�H��͉nQKuB3ex/�ǖ��ӜL-֭�R�ײ��#R=c��^�ƺ����`� �$�$M�h[�7��_<}tU���D�6'+uD㱲������X&�5>�g��hVG�f�t��u��L}�����Y��&�3Gc���V���k3�Ҳ��͕�@�nD³N� ��C�l�Q�#�Ik1Q�
���8�l�bFPG�@��PB*|P�e��@/��L����Q�k0�'�m�&��l��6�|h�t���q{�'�h���8�(�y��w��Kq~ٵ/�̧]p%=�f��[˸�*��[�ʜؿ6⌅�*����[����G@�b�@��<��&�݋�]a|2XBP�j4�u	mf\���5����7㉀6�:rE9c�q��w*6��a��J�}y�j�Ə��� �����Lr�g����k��sShQ;�`�$��H����AT2F�k1�"W��XS,� ��%��B43
��Ҩ�Q�%�&s}xp ��g���JqQ�1�d$��k�,a�ː�n�+D'�fTj�[�'3Y*����'A��.��2��e��f�Ew����H|�Oi_�e��&��N���D�1�q=Ǝ��MF�.�-u�il!����I�.[�.�4˪�i�s�`f�"1AX1�3�S��p��"v!�څ����.i$w����*�?�Թ��9;
y?��(ؼ�i�^�(�R�!�e"�ɸ)��|�it����J1^c-C5_,���9s�����S�k��������q�,�'���a)��q�;����~���;�a�;�[��d_L�$ �Vi���C5����Fҭu_�:��]�.�"N��,:�-�>��]�����$�ɿ��m�[�bx�ol,I���Uf/`�e֣��dCPr#�';�V��6p�;�p�gy�ݬ+a�;]��]T�Ƹ�ʿ���V_��BA�,�`���&�O�K���De��s�u��0��X�!T찥d߲��	&wMI���Ё��~��"��4j�q d����tbi�El ��D���`��uEW�K�R�wd�7�9�c�"�U�h	+$������'��J�V#�b�W�K��(y�	����R�e���kڎm,�(^��ȼ�=�;�=uo6���yQ�$O�6�{e���%(������/�q�2��ρ��T�r�}�=Z~O����������_��d:Y*WeAi:U��F'N�ݭx$ଳ���|M�9�Ed���Y��6����eI�o�5���M�1�V��N�4)��� �O��,�0��QA�����aH'���*TBʹ���^��ݸd�I���A���]�!�.����>����Tf���(:�g�w6t�t��$��|7@[�g��Q��n�f�D�y���B�B���+��%�(`�h\��\O_Fv�?7���Y1�!M�"�/Ȝr�2l���`�tk��2t\U�_3E�cs�1�Ă��/b��;�Y�HQ�R��c��%Q�͓0R�h2�=b�qD��M�PO���9N���j0��.[����ٿ�Z'U�se��p�Ha�6ut��F��ğQ�.A%NCn�Z�?`^�FF�Ӹ}A�_�+͋��}}"�$�Cu�\4dx�	3Q�G��ۯw��u"� �"�nz�``;�[��3y��e3�x�B�V�gS��N�1�֘D�:c��ǰO��Hn�������`�	p�a�;����[S����n�<��3��9r��#^��hqgZ뽰<:��΢7���B��3Kp�0����4��3_�f=�b�
��a/W��r,��[�A>���$�NP|YW�7����5E2U��;����m�@����ʉ��c_#]����'RK�a�4����,��X�;��R��~#���;����㪢Dt8�KS�{��U��oU^��
c�7�"yjd*S��=�i+�LJv���Dt�������-��">70ߟ����|y�(���ĝ���ėx�R5)�i�8�2��ղ 9x��P�AC��V��k�چm��4Vt�""Y�$G'D}-��n��?�z��`����߉��O�'{W�)\���E�q�h���Z,/��|�M�*K}b�mխc��+]�j�t-�IN ���^J�9�Ӏ�QBWY�R��<�oQ��"0O;1ؼ%�`m}+l���s�װ[
���^ȱ���qu�Px���!�.�W\s|����:4�`�z[���$�Em�����ñ��rfġ��I�_����FWI��}+*w�|;������ٲZA��sMb�Pu� �T�����j���b?xI1��:��yCֿ���Ô��n��k����N<���.U?<^�@�7z�X,��"�)�!d�;��(rlz���4��ɕj���J�Pɀ8z!��?o;���n�` �	��Qc�{��P�q�d����lA����Ο�(����jJ+��텖g˂Łؼ*}������|��$̩�V�V�(+e�����E�*y5FE�t�hв��B��`{�����pP�ghD�h�P�7���@ޫ�(��T�6�����1�� 8�ẇ�A:���0�%�� ^����ڏG��T�4�Eބ��%�����:KDݜh��nk'CAh	
4:졞[!�Eϸ���Ǩ;�~���
(�b��e�nT�EXl�t�/2z�p�2x�I��b�����g���,M����'��$�vu6�f��!�� OQ�D?I{�Z!+��/G6~�ȸ�74B� �TX�'�]|��I��G�@�n�q2�������^˟8Ci[C�1�!~�2��c���������l�@�w��l�;�U��"��w�k͟;����d��O5�eT஢��҉`�V�W�e6j�"I�?M[�i�!gT+%�NiM>zI ߪi�}�䃒��s�`�	R7|���&��ʲ�ySA��>9/<k��+�F�`��V,4�H �Χ���" E��Qpwdy�T�I�[�����XQ�B�+��2����O�@����>+���1f�1�T�H�Zo�p��)�I�)��c�~�g�z Q�g�h�tn��H��E.R����0�y�R���d���4yȩ_�{�Ws�g�1«p��;CI<2��C �yKd������\�Dnu��F�֡K����A��8���~ 5������$���邑�Lh� ��z/b�[���U��^����dh�}�b=K�/�K�*�sS�A�r*
c����t�RR�$0�螷 	��Q�+=T�EC�q["�=�`�:xV��d�@�}����h`
�2��i#B}�V���:Rc��cLr��1f�4��47����/�5Kf�}~�G��xz')�;DNn���<�sV̙�kىi���bt���P%�)~�ҙ�؀ы+���h�5� Ǔ�7Wb}ߩ��J|}P��s>,=S)�
�x~�	�إP$TR��W�6ֺV�8a�*Q!�ܥ�_��3�����F[��L�'p�(]��' �r���D ���>�Br�[B����G���>>�{��'��0+	�w��Gݨ�F��l��!�0Dm
-����2!� \ \����V�G�|����b�!?��!��n?�ub/��˒
�[�c�`wc�z-��a�lq��6L-�����k}��87RYMla�g��"�C�qn��������u��=�	�K��!�*�#��!:8{"m9�K�{Ł��/�e��G�1T��V�,Zg扁<��������n3�
뫯-���oF�h}�^*|����&��NXѾ�Y)�CF�� J���-B�Oy�5���h�E0
k�����i?h�]h�y��"��K)�&}�|�Ȑ�Y��{�"U�;� .c��3�������g��3�E>Y����x���-��I���U�\��	GN3�ZY=sTE��ε���'�Ň�-DR�\^K��/s�F��d�g�y�.ѲF�4��}U�{F�QNK� Asn�rP�%m��� #�x��_�t�G38�@(7si�#5@���M�8w0D�#�����cS�O�Z����V�-��Nφ�<�)d��ب��T�����Mc|�A:8>cYNL�7Ň���=�0%���V�O;4QO�3�p��s��g�&�A�����v4
��U�z��	�\��(���藴��i�ia�9�̙�3����~5>?:ڲXD�#gA>\�jͤ��=�[E����F$f;b��8��y��5�1�UL	S�`���*��N;F5#�=�0PW�v��LOZ�Y	��y.Z��i�Im��GM'�Mq�ºS].�u"�+�C2��A[��0:+7A�8Z�v������zw�v5��F��ku4�L���"��.�0���ي�L�z�mB��=&�)-�t0�G��>���B����j����a��z��_�=�R3S��>^:5%�>��p�A��� *�����;'T�Tz�m����A�4R�,Eg0 ��GK��Y��M�|�lO�\��?�K�w��(AM'��0����}���Y�uZ�!7M�h8���I��j 5�d���
�r��d�_=!�~�%�'I=��\v�Ғ�>O�j87C����7Ѿ:̪M�������Ƴ�Ǝ����17�R��\���ܕ�ɐ���J� �����DY#���J9�f���Hiǖܸ~��%
s�0{�&:H`��/���4;�]'��F���|�6Hb�Cr�:^!$v=;�c�H(9p4M��_���I�R��>�"V�QUp_
�n����)�lіi���0�W\W��B`��x���	%A��T�����id-qm��e�qx�b�8�ܘ�?U�0�/��_B;� �"0�./\Cu�P�M|��_��%?n�S�|�Gc
2?�$5a��Yh��X�D�2�8���߲fTǦ�l26z!���g<is�T[}#��Ũ��%��8����K�R;���̞d����
���p��&؃I%����JH�.M�AQ	i�3������{2���(���߽F̳S��PKa��g��ȮAg���3�����S����+#�ԛ�����q\	5���%P��Q&��u�y[��Ak����<���B��=ڽW�,�=3�`�[��=��%�߷_$kS����B\���|ko=�r�Y���ʜ�P�_�|v�>���kpF/9�|��b��q�)Q�+��Ig����*ݿ����L۠\�&mԎ� �ݎ)@���� �X�2:n��P�C���Z8̍��A������ӓ  �j�a"z�li��W'�H["�i/پӤ�h&��	��
�,�fK!ͭL05�3����-�A�9X�[��(������,X��3��来��!�_D��AG�ĳ~?�-�h*����wG՚A�h$Q�zt˥�'�u"y��u5fo]/��Zl�	����1�GSCP�f�mŵ����qJ9�@��H<\���$E�T���=d�+[��6YݵA����2I+D|�s�q��TO{zE�G��?w�S�ވ� *k58S�d�B��&Q����n$h@+z��|�)��	(\����LX,�⸞��c�7��ђ��OU�R���sf����Fg��s�o���>�H���ȹ�����ԳEa|$���R����Q��h*Oxa,1-��b�����b�K��UB�5�l���L) ��uL��6���w����P�^�h��BL���8F�M�[a����&W�G��+&j�&�-""��%l����o��k'`��_:F|7أ8���rK~��fQ{'u�_i(,�@��ϯbE�P��I�-�0)�V���F�]�O�!4M� ������t%D��FW
9:Ց^�HL�f'Yl�<����!���$S-�eJ+��q+I��}��NoVZ�
7p��j��g�/�Z��%ֹ�q*!�Ӊ��ϒZ?-E&�sH�m�!,M�+T,4�y�!@x���w �p`I+�	,xx:�5��ȷ�l��2a7%��8Ȟ6�i���
�g�4�6Y'�e��>���P��$�ۨ:L�0�w�`s`'}NW��*
�@�'�D�ӡ�y$P��r����?Y-�O�6�9:z � R�(rՒd��P��	�2�$H�*Dɂ-� ����	(��6V��WAa�|��ޑL��Z�J��E����J�M������:�YK\\�����ha5�ry�y�4P�&͛������eS �}JqtG1�4�|`�� QG��&fa$?B\}��o���,,��S��^`Į�hy�����W����=���j"�Yu72�����H��d�Z��f��)7�L�Gi$���3:����ݙ|U��G΍�����ϫ�P �(�)I��iI����iừ��S��T��~~C�;�z �&�Ͳ��)�KE��Z�+���jcђ`�C���ʗA+�]��Dh~HlZWM�z�_xXo:��(E:�!�- �q,�����da
���Zz�`x�n��� ART<0��c����P��U���p<�X��ި0i�|E�� ��K�6�h8�a��̂ �����$BY>��xs�mv�T�Zz������4"Ń*�����@-H�	��s�	T8c�D�F��6�d�n�w�E|*,�8�,R�r�z�=b[ƺ��#�M�ꊣ�� 壹7Y/T�����g�&i~��@��î��fX� ����~у�r\�5vZ���?jS��j��B��>6�T��/�!p.4�ؚ�K�D���K{a��ן.��@e�=�*8��������>ux���k�� ��L�����>D*��ʒr�,�z�=;��m��{4�i��o|�k�?�,����"�t�2S�O�^c��>��pG���&Z�	U>�Ga/��z�4������R�����$n��a�}�t�����RN9�f�K�v���Ui�K8�F�΋���3\�O�7����.,�2�(߁p��n3�~H	:8��)"�y^e@^7���z�1�=&E���5���)�#��&b�-�FiC�;��l`M���T�*����;�oO2��A��=sIwZ~� I�[{@��Q�u(���6dNnTZ����Yk��`���ո�J���/B~��<��6���P�1Q��ljm*����FL� 3���yǌsnG�r�/,D��u�V�p��h�:�K�S��;�M�"���P����%9j_z�#��ȯ�'�Jm�N���L�?��,(x�<:��ߜΞW������'���L_>�E���"ZeIZ�"�c��>L��N�MQx�>K�4  �Q/΋l�͐����U��3��*̉�3�"%!�šm�â��;����=�j�,̖N�{���zs�_�Do��1!�ڂ65v�ݝE����xRc�K��JaM
ő��=-��!��S��`���u�W�/�ʱ6Ӹ��U���t�r��Y��WT����U�	a�����Ug�o��ؙ�;~t�C'�����[�������=�`�\��r���Q���d�T0��+�e�Qb�c�J�()�����A2 �)S�RD�L_1��~'�h�Ɣ�Z���j�QN���4@��4���b��^s'܃�f4����7�A��3$ r�G�h,��e(��{�h���w>V��V��(B�zF�EV7|�P�J��ʱ5#f��@/�p�N��gg}�L�zM�����7U'�䋜��y-��ny�<_zbj0PI���K��Dk�x�:��r�J���r@�4S/�&W�{� �"zda��jE��]Mg.;�_��G��e�v��?5�iMB��IP�'�_*<�xJ$���cQ��.G#�L+j8Pvz��Q�覝�&�CI�.P�/h5>�T;Pi&٥�.c2	�Z��3�h���.]T�u����ɧ��!��j����p�_�������5�Rn�j�b�]*T�%�.~r��v��%�r���O'T��9�U�r���=��QX�J������Fs������q�U�VUS-EmqȿA�MJ�3��#
i�R��FAޑG�y��.��r��6�X!S�L����h�=w4���)p�6œ���|A1����64��7X�Ҫ�T�8�Xl�<��<H;r���9p�c��>;�����|JQP���m�Iz��usWq�b[�f�;E�Pä-�]p���:�v�mڦ�v��SdҠ�J���W.d�����D�u1�o|ñ4/!�I��}2�i�����wC�w���#�Ϯ?,Ц��Uk��16[n���d�}SV����g�X��9p�/��[�����=c���W,u�X��Ո���f,�/��w�Ɣ�̯�3�U�xjZ��䮣�����h�a�����k��+b�v�ɫ��(�Og�5�743p��nt�	[^L���ɩu�����,�AL�D�ܜ&�w��Vy���)n��s}t�Ѥ�3+U5z1-]P�5��a��ķjO��q��o���k�bf,z\�#�s����!h��6%+�lC��d������+u&R�]���+�z�t��u�^CǑKV�]"p�����1�Uk/e�������i�پ���M��D��M�����1���F��E�B�����=<wA���	x�!�:�>fUGޥ:(�\�`���	r������G2m��͝��u�'�(�����M,��X#t��@5�>K�M��E�!8����̏?w�ś(�"��^��N��������T��\������Z��J��c@fqdi���(���_���̐hJ�M�x����YU*0ȍ7�rE��;ƾl��в���j4	�����!�vg�T�x�sP���
@C�i����7�J��t��!�8���,�w���Qס� E|g��<��+���U��0+��t"5����k}�����A&�!P#k\�ƙ���R�1���E�8K^J�#�5f:���`E�~{�ѧ*	.I8���ʹD�p��|kU}{
�%,��R���h�#Z���L�1	.�Ǭ^�,]��B*5��t�,/�t��a}N�,˭��NK=��|o�ʿP�:CRF6��jT�2[c�4���A�G�r���q�g9��el����c���}����G
 	�w�Շ�uw/O��g��<&��cy�����O������� ���F��+�4�
~�6"��=\9��r�9ifA��sJF�G���+#���&5ii��yB6c^�k�n�%q�F��&ʻs�G�]9���ӕ�����ڃϖ
R��j*���|���g�C?��{�6��p��Hɽ�Q wT�X�-%��l�@�1��H�s�2��ūd���QUaX���\��shh��G��g��< ���jG�8������c��V�D�;����=�^F�~S]>թ������%l�[��G���&��E@�jeK����/Ȯ�U��#7~�@�nI:-
��O��.e�m��Z�1�W��vo���p�̐��ډ��������׽`�.��u���xR�v���������+O5���?�,s��{�]�����q��F�F���ZJ�43�T	���0�NT�u�}�p_V�K�Y!16�Wl?�W��*�9T�优Hhq��u2̅A�|PM�'[� ���	ҙ������c�^�����; �l�ܸЗxU�JkM�_��pkq��0jk���~%�f�璡��g+�	��yF�c�rJH4���g�H��Z�Pm˛
�(���M6ɹ߫�J�^�!G�yt��@��Ǳ���$�����;a�P�F�����WȊ�g�r�j[���8���,��Џ@顄��no�cX�'#�R�>���;�\ְ��AC5�R6~��N^|1�*������{ "r�-vy<rK��x��N��C���A�h�mM	�ā�}����48��qɫw��E/Qnr*�[N-q/A�N|K��ac����YV����ӿ��� %}i��A����mGRgg��D��&#
3��U�$o�	;D'e��%�u�JL|����FC��ezâ��Ȍ(+��r9h5�D�ks��8,E��t�n�H�a�)�7^9�H�V,�+ڳ��\����шs�?]zf�{[���5�C�~�5��Zi!b��p�#�
]��q)XJs#�u��L�fmh���"�yi4�a ��(8g�`c��W�F�f&@
���A!Mq����1�wy-v�˘�4����d�l�82��`�x.��HlXultm���<o�H�&2]Q✺�*�8���:*����_c��	_
	.��罀����ʽ�-J�Ȥz|O���| k����zxcu�<;H�2-������Z*g���E6�%�hv{w0����Ш5�1���xy,�j��a�)�7}���]l��8*�Qʴ�f'�W̃��A͚x���?�vWR�^B]D�yAЅ)?E�9!��26�ہw���)%�6�ZI���M�K���9]�"�m_��L
41��DW���c�ѽE}��h;o���:UW�|y,jɝ=YC���]8��p����S�~z�PU�.|�� �nT�o�V`/-��L J���nN1o6@WV>d�L�i 4�?�?dWf�k/l�w~z���4��A��/]��v��~���&F���=s�I��Q�<x���UaR	��R�Ī����F��(F�ћ�Vt2��{�Z=��{[��VB�`���"�i�EN����\�j���;�`%��l����*ey���x�lCn��zk�\��aSWG�2\�[�W��NN�I t@�~
.c�����xT5*u�2��b㽛x�@��(ޏ��%���4~�y-����ѱ�Hw����a%��Qb�f�15�a�F�Rn⭿������"򙠓ee4�O%%���.k��|9�شE�OT������*+	d�n���2h\T��0|,��Wev@J�g�y���|�y�y��c�}ץ�i�㠩�t:"��Cq�)4/�U�l!z!�Q�0��kgY�3��R�<���^���Dj���5'�@��!���ɼ�i�eͨS��q��9��#�É��@o��&�ǧ��d٠��$2m��
��6�)�Ŷ5C�{��Pǝ�|�>?j�_罫z/��o�Qf>��
�'�Ν�c��:�|6������?b4K�[�M���k�'�^Gb��B��O�����?�kv�B����_owN�%��n����=y�d"��#�2``��Md#A�H����yWW�_LR�qi����y}R�M���{����]�����z`�/�Qw��،��sH@�t�L�o[�r��i���$7���E�5+3����#�,6@����B� /�lH�M���bn���a���#�\������B��¿6J���><�' ��tj���7�j
�D)!��f|ד���?(� Ä́l~?K�iX���:c����kR"l�rʐkgv���on��71��`�?�F��K����3��S��ջ!�,̱�9l1F�ԕ=:o�2EFi�8���Y��
Of�҄.)*�R��%i}��C�\i��0�i���t��$��E}�z�Do����`]�;�t�>%��bOҶٻ�e�������`�3�($4�IJqlr��������v]k���P��������l����[�� �5:^�#e^d��XVgQ���G�/���9-��o06@o���������	�ҹfF��쁞�D|����������K���H�W����ք�@�#�s׌�4��0�?�]TA�6gu�-��{��WBNpl������a:��X~S�+;��KS�hjȧL3 g7�
I|ͭ���'o'�̜[�٘�<8z�&%ϑ����6&��-'�L��V���^��rf����_M1oԔ��A릇�[��C�����$�������9ĩujh�AY(��G0��_�LS���W��?-�r7�o��8b�G�Q�y	$#�����K8�'�|�4�����4���������>/;N�Y�'ļ˅*�0D�i���'���S��	
�qQB|�o��&�7��Y"�S1�M��L��Ծ+�.!��>-V��
���o��{?K�����Ÿ1f^�,�����͵f�u�RW�����N���;��k�w�CC��E	���t��J<%�����G���\{��y�+���*�p/��4��d.�D�c�6Pʜ��un�X�#�=�P��d�)�bJ�nT0�-��)ֽ>'��j
5�����P1�ٟld�����28�u�~*��"�g���*�$R}1�̗���g�l�T�eG��Z1�J���
¤$��lkj��=���'	x���������9L��9��O�F�����y,����4Z-RUC���;j8�|7�����P����Hw�C\ ������|�z��0��վ��k������"�鲡�d�q�ZDO�(Y����F�D �Ġ���hQB�Hj���QFA��R��i�y�ܨ�4����
0P��<K�z*!�����c���RT��I���_�Q�M"��B��&$%#��(��Y������p�/%����e��u��6�5��΁�:��̇��>$�x�uX+�qU-T&�l��nt�C���Rx�>�2�����͒)B<$����A&�w����y6v;j]N� ���c6ۚUP"JVB-/��3�R��;?����J�R��y�|��] n���$�_ж
�X;~)!���@ _[��[=<�V2�0q�קŕ����0���s�N�՛�S�}��;vQ�UZ��ŀ,����Yq/C4�����n�9 3�p ��|������җ�{��#�"���J�r�Q!�D��+�zkg�h�����Ky��1v<��}� T�D�L9�������D	�d;�k��S��5ll*�����t� `Y�9	�����WA�*U	f�q|��X���I9�'���.ǐ������b#���HZHK���
6�Gk��1<͇�"b"O�l߲k�Ȼys������;�5G���?���ޠ���-��Y򻶍����J��&����j�f=,�����-�G�o>�����/�i5��W|��)���T>qf��,3F������Y�����
��ZY�͚/l���!�V�G����UyR��%�V�B��Y���;ޣ#�^�C��ֻ����-�F�����*���"@��blu�\ګܓҋD�B��p�h�۷���~�P�+��렍�X�R���X7�e@���,R	�sؼ�P�@�2L���g�_�W��Q����4�+<��ǡ������=��4����,��O
����>g���ɿ��%����"Э�f�w�e�+����`P~��O|n�Dl�^y��/Vv^l0�^����`ˢ9�WL�LQ�y8�o g�`!�h�s�|{AP�W�OcD�14�oԹ=��N4��,o!���UF�U�dB��"9�s��$a�1��{�G���2��n�Q�;s�]޻�S��ǫ�ƕ:ڸ|��<�
��d�t!�%�o@I_�B�5?i;������ԅ�2�0?��Y��5�Y��%����@��!oܑ��/��H�*���]F���p�t1n��h$� ʶ�o2:ޭD�L��#�f��1��L�@�' ��H�0�;)b�@�|��%���:�܋x��I��j�+�׹�Ԝʰs2)�,�30P�䫴�T���_����'���fY
S.nj�Q�TC���©����QX0C�z���>w;�q`�W����d������t���vsŕ{_peq��,ht���E��y�h�(�f�Į�ċ7:!��@�>�)���+X'$��#O����l�x�J�7��'G�~��ٹ[Ə!E��S�����%�+
+�E�2�����U�~倬n|'�9Z�P���eݰJx">����C�B1��vn�B
����Q�=�+��ؕ1�mr��6W$��zE�6JŲ�ͦA"�A�˴�^���6�[Q$�$
��#�|��9v�*KΡc���>�6w8<��}Z��^��h��S`�"jp�g��J�$�^g�`7��G�s�y���1��Yj��?�w�n�.&�����&�c�}X�c�
X+8�D�'���߫b�st��Xs�#'���v�hG9��c-[���ջ��q����O�&%)*���~�"M�u�����x����A���W]��`N~���|xr_�b_;s�P�=rb6ϓ�:˕�7���Dϐ��(^�gf�J��=nd%�h�Mů�t���)�g5��\Pi5l�Of��ߣf|2v#!������$���ܪ8���땍�/KI�(�tQȕ���_?�, 哪U�c%'h�:.s�O��C˵zb=l)tp	]�������<oq\Ѹ��5�\���S��m��g0pޒls[>��=�_�Q�*�j���-V����Q���h�İ����g��r��𒇫X55�[����O�I8��z��՗���4p��9cڞ`���ԉ��_�������v_t���}����#-���6�e3�Ǒq��ˊ���d����^���qܧ��z	��mB���YZ��jc��1��m���Uhg����4�}A�Q<�Mg�uA"��t�M��5�:�1Z�}�
�_��l�k���)��˃,���?�x�1�:��>�]1��&MSυ�Y�W�EƧ�̢)�<�LA~�v�P���9*��dU�mP[~�\ul{�ƴ^�E���~��e����@#ϰ\��:0�C��=��Ж�O�Ys�I9���%_����Y�>�͞s��A�\�J#؏��IO��+�z�"��CedF����}~8�T=ݢ>�D�cw���}�1PT�Y���RT�P��$���,+�mBg@hU�x1��r%Fd��%b�ݝ�w��ؘ�mn�Y.�Մ��A�}m��VԾ��#d=���J�'���8�w����X��}�;��<�;�����π��AJKdi���(���@�?ի2�H�� ׹�ҷ[��9(x4g��w��5��0�!:���Vt��=�
8ӥ]��SЎW��N�Y�T��m`��hk*���v����T } Yo�����?��o��y�Pƻј:ڟ�OHe��c]2*M�/]�����`,Ǜ��`�;#A�L'I:�,,5���7�Df��y˱�6P6Ӿ����-9�-L6P>��J2B�d�	WvџJ�����v6�s���ʝ$�?��6"9��Óq��ǆ=�x�?��7�d�b�+�y��s������~��� ���7�-Y�&��#��x=!(��,��O5�����9P�8��!3�0FP��[ ?}y���[�t�`�&��\�5d��n;���5�P9L�|�_���0dEn��Ti�j�$\����uc�9�;�_@�3~���H$X=�ы�����3�®�QA���'�N��i��@�x�Q��k����p?P۸��VJ+*P�ѥ��\?!��"�%�� �Йk������t���
�&�5���#ew
���#l�g�yѠ�:!|u���nSz��`C��)�_��{
�N&Wm*�#)��['��.��TO�L�:�D(��jZ#����l���Al/���DI��G�U�8�� �͚���М:���+\�EƝ-�	"�]�44s/L����5@�o+�Cd�#��q�l���=�տ�E~0pQ���>�`�US��_��R�t�~������������ٷ)�Cj��kHӞrbU�f�E�SP�#\2����&��Z��xw�M�/��(9�4�8	�R7�G��$��E����l�Bk�[9�%�,�G��>��y+m@����~R�p9�W?�`�!5�U_�I3H0���OXkfU'�1!���_V������bH|Z#]�(��F-�0������_LE0��5S��a(&�����ڷ�؟`ؐ�cN:��t���|�~C�D$�'� ���7|'���7��̼���m���n@��[-n�VݽF%l�]�X���� ��4���M����D�Ɗ�.���}�s��ﺑ��=��;xꕐ�şhu@��↢���-�K�ON
���v V �%YQ�5�g���~̛a֜B��Zq�ƾ|��g�ߍ��K�+�q={5�Ц{�N��m����n��M ��b(��+�[�%m�7w&�3=J �����	|W�'r�P��a�i��ؘkM2���H�GJ�.Х஼2U�~�k��F�B������#�7�~�ID$��)(VBS�Ř��`�N�/GQ�:;j.�D�7+�M����8����ݼ�+�}M��rR���Ii�(���g@C\@Q8ci�.��Y�3�&�R��y�~����p��%a�� �
	U����X�,8�ԊF,CE*��i�'F�18�)�Yo�D�^�1�Ԋ� -R�xG4�SP�����,��~�J�1z9om�dR�V�Y܆��6�!�K8
v� n���{���RZW"�y����S��h��H�0�r9��<�<Cc�H�n̧�De���;�gүn�g�M�M1���ּ3gIY�z,�Y�n���l�3j���|͵)�Pn�*��V=,���-S��0k�+G{�J�V�� S�^e���������b��PȆs�h�K{z��X�*��
^�%�y��Zis���fR���x�{Cɡ�����1�5�Lu+���Yi���jyq��ծV �;�3�T�FK�y2������q۔.��Mi '����s9ﰐ�'���h�� �9�i�M�o!��̼���_,�eSo�[ ��z�E�/j�ZT9����I�Ÿ�wrfkP=vXA�{D�?=Qm���)�k �	�S�ԉW�Ն��OU!:G��0��v�}ן�9-���H�:���`���ԌbN떖bd)��XW]��8 �=}]
X�4�e�v���VG��x��f��������#Mo�ꉏ�ȁ��/�D�LrrV�:�MN!����qK�B1�H��f���J�x�ס+BjHB(|�W�}hi���spJ���@BL��0v�vH)yXV�sm���.'́Sq_�Uo3V�.(�x�ݫ91���CA<�훩y*�~�Q��d�uo\,��
�L� ��yL3&�@k�Z�;|��u�?�3���s#H"�w�W�ٹ����.G���os.8�y���d�Mn>�+���V�(mD��'h��2�8����Z�s'�n��W��	����j1BK�t�v�,�������N��A�k�k��E%�����4"����$�x*8�@��� '�P���7�ϼ����pLU�ġ̃����樤X��M�	 6z���f���/!+e����se8|�ꂷT��|]o?L�l>6H�k���
f.0�T��mI���"3z��!��P�$�JA�M&;�Z�Z�5�KVK�tK7oD�ϩC��&��4b�������X_�0�"�Z{x�}�{�d;x����3+{(ۧų�WJ[o_��i�7ᄄfV[�U�y�β�d�h����nҼL��u�H��8���^DlK	_?���h@�#�h�^���k0�򌻣��H��2���&^�M��s;�����.�^�21iͯ@����ΰjC���N�m�����[;��]
Uc�"	�����4=��<�wp����R�,����k��Y4c��_3Z��W����ru@������h{cz�?! ��s�{��ɳ��=��Yb
�J��7��$$?<Fs"��&�k��}�AQ�s��� �I�Po�{�+5��٥�C[I��!�����Mk� i��)Vه��b��bm�����h ������q7uB+�$�ઔq�瞣� �����:�U$������(#u�N���]��{~��3D�;�L��g�{e?��d?�M��X%dD���*�`��� �n��������e�Z��lU���muP�MDa�w�5d���.Y����`u�R�}�(w�Q��ѿ��o;��6Z4ѵ��^���P�!�_S�ᬅ�ؼ�)F�A�^WD{.ޥbyu\���.�8�G��F�[��7��+�	WH������%�&��G�ʳ�G/�UI3�ry^�x���no��o2-�.
�y,���e��_�g^����WH��D�r��Z��<i:�gٗ���<j��Qt@L����k@ܫ�N���K�s!237c$��B��>Qfi�9�3�P�F�u�9h�i�OiP%�#2��x)M��ϙ�1}���G3�o2��S1��;8�NȖsї�[[�H"_�S�%���V,�C�m.�2�{ mW�R$��s5͉�8��#(�\��C�r�d4�k�}��������h�������D��i��wrh]�YQ��}倠���Z��id�h�&�v�x�Q��U�d�S�f���}4����5�Iyo���&%���|���8����/�o�q�T�j]��sؘ�������4��m�Ցt�i�L��`87��2v_���%S�1���90�6�y7B�ԶZ�n����C�h�nq%�jiM��\�wR�U���>���+��fͼb]�X�n߻?��f�ن�����O����ӕ��0^�{���Q&�"8�5Z7�e	��fW;r	���:'!!�J+�UcԘ�Riŭ�#�˨�'����j�(b��
����kM	AD�Y��!ɀ�T9|ۑ�a���g�����GU�S=�ʥ��k/��d��*�d���5��N�zLX�����Ж����	p�JzS���*�@N��2��t⭿��y�">��4�����F�fܶ�>�E����Yp�y��<[7G�τ�T0�d�ve��K�\��4ma���D�V�Y�U�EK�Y�M�pϰd��J�e٤�K����V�g���SX�P��ǻK��e#�K��i�=�G���m�PO�.�����%K���jI�|k���	3Ot$c�S�_��y��l�x�y�΅?RZ�����N�[ ��)��� Sg) ���U�.�% �>��S�`ft�r%��� R5��M_�F���^9R'n��K���ȫii��e�9�X|0^�v�w�W��w��oz�F��C�|e�B��%�D�d�{�F8���n�vs���Wb�|��Jb(n�BB�DФ�8�-�LQy5¦����	rR��~g�""Rצj����_7(Ӳ���h�g�TN"K��������䎥������)h)��B�檬�����z�];?�Q�K��H�^{[E����X���L�!G�_1#��4�Ad��ꯆ�9��=�!s��77���l�Xw\����B��*����go�&�4�@:�%���@ʔ/{_��{�y_��i����=]5���tiC}-9�)��*VZ�Q-N��e��-�7̞�*H�`P��ԦXbqK#.��:O�[΢8�&���	�{#�׎%��S��r�@W�~�j�F+[�GC_T0��k�㎳����}�5��,دAP�2f�	�u�I��kZT�z���H�3���s6fA�_��h��$�7R��A������>�^�	��|�;�iv:ʅ�k-r��r�:�G�x��h�i�SD{���Ú�xL�@���|�'�-�ø�@�ap��mt]&!DB��z�2G~3��V�Vl�5(��{���8ż �ySCT?�Z�GZ=[���d����ww��Mٗ>? Bzw�����1����tgA�& y+ �e��܆���A�d?E�)N��6 ���\���{����B�d������` h���`U�!xfU���I�<~o:�%�x"ǿB��|^��Y+.{ґ&-������(�Q ����d��"��`�
6�uc������C��DP�[��oʁ���ƾ�g`�*������]�/E����
�����D!��jUةU�8�e^){�Db��n�4l����ƕ�Qwj��Usu���������^��.q�� �i�izS��#�!�c��Qƾ���ZO�(|#M�Zt�%
�<h�ˎ�p��H˾�1�9��NVK'!#0�ϕu	�1���x.j}�j�x�X4�곟�ŵ3̲$�"	��U//Q_P'EK��F��E��OL����dRhF(\[�P�/�ɓ�s"w��$�eqs�<��76��N17��8��?�ʁ:Wi�5�	�u$;p��UH�@����6~��>��BKpXNZQ[\�B�A4?+�?�)��%���F��=M�Yd�u��k"��F/e�
��I#�^I��d�쌁��xp��Ȑ{0�/�0fB��~S����s5Aq���]�r�倨��E���`\*��͂d�qe�bTI�xRzU �Ѥ-#��CT$�BUۃ�a������\S���΄Tt܇����c%���	�=�PV�቏D;p���U���!y|&�0�F>O���,�3.���k�"#]�^wM���2��9PK-	=�֐-{C�-,STb���DFe),��`�1�].��ʽV$���P�7:�eRT�`e��ӥUK�pܝ83��6�p s��N�(�~^�c���%G��¥ŗ<�3��р�����>a��x�!���y��md�%��΍���=������2��g���PR�c��Q�-o7�j��$�1F<_-N�-ӝK�渦����t�|4\_�eG��b6;ޑ�r3��+��v[4��.`���l�K0I�*`fdp�S�4�}��]���A8����{�P0 _�)!��˨��$į�<j�{rcL�v����~�00��$�(Ɏa��T������nixQG�amD�=D�b�B��
�������]Y�X��&�\�5�w�=��()g���E:���,ُ
�#O'�o}�D�Q�ȱ�-�ĩ��5G&�>c$��o�5�jV�  Tx�i!�l�P��*tЪ�iI������;V���H�J!!��i6b��LW)7[\](�E���Y��� ����	��u$�f�qn�
���8T�!8�`̝�]ځ�b6yJ�?*�5�I�)\"�v�=ā^��X�t�j84�K��X̟b�� T@�+���,'�S��9�}8�`��
F��7D`�2�\��.΄G�uR6KP �%�L"`�e���a�p�[��z�y�"�h�l��%�g�>��x`�rY��7v��1f�b�0&i�H>M��+��.Z��u�G�'d��n����՗Q�ԟ{���V-�;���mh���1�s־�#�L|��$=%���Y�H�j�Q#�ύ���%sme��Y��Z4L0Q�EA\���C�>�M0�<3*]���,pS�G9y��������j�s��D�D���֗���jG4�Y��\���vW(��(Mt�qG��:��l��m�R�{H�ͺ�F�}�O�c���x��W�Qt�+܍��3�sEq��b��5؝ibD��W�-��x97� P*�Â��ЙC��}��;�}X��V�|�:`L�H~���Y:��n�x�W�S��k�s�:��]��P���9@���ʿ�M�e��,���B=�S�2�1��IC:� �ɰ�IPʴ��Bw���Í�dj�&'��9!�?���(�o8�	��zN!�8w�D|��9� �Oy&\�ʨƻ�d7=�Yz�Ϋm)���&2�4$�qn�G�^��&p�P�vau�9��*�+\{`-��<'�͎?����I�\y�ȇ8���"y>x:����)�x�hb�ɡ^�J�ݬ�s���޶[��Is���Hp���*�����]A9 <Er\h|�H�A����oB��@�t�Bw˰�[G���kaw���h��[����Yn���U�X-�k�K��H��C���QUז���0a%-��x��*�u�I�)������+�;�Mgڏ�Z3���75�ntObG6�ݮ���g%B�BF7�Z���d��)���n���B��Y�nU�Ea�^>�ec�D��н�+6�e��yh�!�0BbSƽ]�lݺt�NȦ��q�g{cXbR���kBP��*�G��s#�#	�r,B ��=��P��Ɉz�����tTZ;{����K��g�V�&�ha_ɼ�s������� \K��L���L�ۮ2�MB�(V�$�F�T�r�K>�:x��
v"����h[�L��m2�Nc�����Ƕ2�{n��˧jS�R�;݋o��:®�9�f2TN8ä���"��_Øm��T?;ن�8����`N.�B���h�I����Zά�-��5�����f�f+�t���|1a�@��Ц���a�ٿ�KA��*�����nTeP�V��ƾ�_[/�4^�� GB�y�珠.,ɛ
�YN\��'��A�����b��iz(�gA�1�.o�^����l��q�a��.J����f_�yT��(�_�d:���pt�菈����2�����d�6|܌*hP�� "���s����2L��p��g��?�ǥ��ULy���2�n�=d��+������.�7�J\9�)A^h^Mh&�*ȁ��g�a�l�ű0NzG8��gF;�:[R�t[�h%�n�͕�.�-T��a��%�!Ba2�#�����~'y�����_�ot��z.�^�
(w�\��`�
9��XG?5��Z�h��zP���z��j�h<�$+�p3�����a�r��^ȏӗ��!���X��=�܎�{i\&�O�m��bg>�Ѷ����<���/��ɰ-C�P1S·�.�?��֝^[je�����\��t��r�^�2��x��+}� ��@�^���t��1����rh�*S�>N��V���<N�����5
�q�!@"��{�M������Q!#��;IMk�|�	�W��^��;5��+�L�9�Y�����?Cy�c�6�tj���������%o�Eyx͋n�n��$,��X�_`�LbH�"�sf���3{�"�U��QX�"�!��sP�(K<<sqQ�����U�x��A��,�܊Ng�&V�۸�\qF�T5�������Q�}��ӣ
Iߒ�����¥"�HI�\pOH�7�ua��^�DC�AWp=�� ����3���p�W�.���VTP�_٢���A�>\��i�;��y��L.y�w���s)ÿ����  ���`kѸı��P���kwu�?�B>�v�J�4��G54����X)lc��6���xY$�Ap�٠hw{(�V伆��#���:X��q%����)of0�����D\3�I6;MZ�z��n���ne�'���2�B7��i�a|2~I)<a=h��vV{��V97��)��3�~Z���E�`,~>����"�	0�X���&�6s�sn�Em�<���&Z��+�K�H��2�P,���#:�x�^��y�Fae�hf��Џ��)�[�)��$���v/�Ր�Ơr�K�qw3,d��^����Zdߴ;����t7�:7���zm>�{?�W�ZMiʢL#5K�Etl)�\��5�g�x6���Qߴ��M{�=��`�mXB�e8��2��D@SkAy�X�v����+I60���/�
��Q95p ���7
��W��A:�_��P,0r� �u|�B������d�����(Yu:����k�.� g��Q�TS���[u����e�͉�.�uRܜOp*X�rg��N�������#���1�Y�c�jf`%`�\��C��Ӑ����x;W0Y�@Yt���ί�� ��?�V�8�bX� �e,�|s�z�fsB���Ee�\[�D�&�iS&*����;-�����W�Z�����%j�tEK�#���U�p��� ����X��t����/x&0j-�a�x��D���oj���3��-?�k0��x���'�=�����$�a�[z����Ŀ��	�:C�n���[��lf�ۈ�� �
�a_�����m��}!�_���#��R&��uv�N0�Wql�2u���H����̈́��K0[���B�/� iBX���φ����1���!�7�6����~�17(���W��BL�1��ξ�2��{(]zo1���#�1��C5]R��m��E'"���'��nt��U�=���}Za�ݛ��G�N�}���	���S��Ě�^��I@^��O��:�̿���W�y�v��>�u�'���d�v�N&�.D�T5��}�D!���N+f<8��gjm0�њ�*��Hę�n��{Wu����h�Z@�3�щ�X��փ�x����Z�� 6�z|U֘]ч���y��]�����v��&Bcʪ�����T~�{ʼW+�y�tl�l�� �_[�O��qp}�^"��;�U[��V\%QJ������5o����)� c�_ ��Z�
(�6Zz~��C���v�5Dk�U��;�=1i��%�bm����gqc�]��p�˂5�NN��{J�a$�#�2���r~6���lG�6�SX���_wu3��0�S�u�a��t�I�t�״y�`u���?꯭��&K�>3��?;�.��3˽ߣ�̀6�X�'b�����XPZ���Q6���q��Ǖ��S2���+��9eL��O�d��}i�xC4A��sC[a�i��	�ZZ�T�
��G�Tz�q؉,��.�8P��(bm.;)k�>�
gR����T�H��
t���U��b��ҡ�s������l��fQ$˵��HuwK�f���m�[�"��S�nl@�P�|`�Q:j
�W�����m,�2�џ!��&�ɮڴ�I�*Pu��.�vv|�Tr���!��#��1�f@�icT��$�����|�s��hdXR.����h�u�5�Ӽ���X�<�U�:ì��yO9r�NLAv�i�P˘�Ar������n��q��iǩ滢l$���pZ9�A}�s �MP�3�vl�+'���	bP��	5q�H�z��j\��p��(��M0vV	�����I�NFm�ƛ�>�u������ċ7�2���c����:��ۺ�V����s�4}���T������X���_��oC�xp�2B"���N�Y��r lEQ��2s�{`or��9[?K��p����g8*�/]����Y
��ߙұ�Lz�X�;>t&���&�L�Ѻ���|R���X�5T��E��`x��;sy��d��&���(���Q��y,��7T���6�_��@�	g�6"��z�F�9����,�~E)|c��ˉt~*���r����O�
@?Ү��$�0�\���T�~�
E��0 ������$�<u`�����͢��J%}�`���  o��� ��rթ�@�D�Kȍƃ)Lh��bي��3��3_/��f6(�a�#��Ir5B1�'F����8nʏ҃J��?��:���!7(�P�NdiS�];}L��ER�"��.��� �xb��e1���LO��V���M�W���֚�/�M5{	�b�#�ș0�B2�p���rƳ����,|"�L��w�����ت/� eR `s��sR5I1S�0i������;�ؚh }�i��8���S/��+����D�ad1���)�V�VXE� W���-���J��7O*������o�BH�}������Z�g ���B��,y}�(
�����%�0�R��^U����Y�V@K�b�ꃽ�`e��Ⱥ�j"r�
c�'w��{���_���_�����E�(�2�� z%���64�5༼�I�WG�Ӕ���L�B�겖�mM��X�j'D��B`eˊ�����#�V�W cQ��>��C����Z��Şݚ��xk��?W����+-����~���~��Y����L�_�X���Ǐ�R��k(����=���q���k�c%@|��Y��u�:!9h|l���τT�be^������@��3�IqD��r���(��NIF�a�v(������`��U�١Xu�Y��K���Q�@b���L��<�����=��:�4p��s3���&��ܮ�ʲ*�?-z��������>���:g���EUǻ��e�-��l���x�q��YD|{��S�f������7f���P����Ho[R��_��A�*@�1��rh���A<�u�(���}[O-��j�)Aż���ÕЋ���i�!��[0�X�r=�v��֓�V3/SU�Ez|��7��A.l
EA�W�����Eժ[�OSѻ�(k)`lt2��w�-����2"^E�bn��rP�f�y/ԱIG���Dy��Ӂ �h�k������Y�a2� ��k`��X���������,̛�-� �S��ao���"kn��cL���{M*³�R��#}п`�C�ƽQ[��>�[�`,�E����;�K���2pm��!M���^���� �kk�e;C��� �?qCz�&�$?���cu�Ss4��
������g��%�}3q��Ɇ����l��e�c��2n�,����͛�`
��&L�������d�jk��+�����2���ΉcO���h�F� 1 �������L�x�o�xkX���)P�p|�ĸ\�r���B%���U/�h+
�7�@f6����݋��6:&7����'�?a�`Ʀ��(%���~DUV�4ԍl�Ju�e�x!�Z��"����vl���ZA�u6��A�">�ښ=]�����5;d��k��f�snZc��3���&ޫ��~&���� g�֣-�r榥l'��Ճ$�%%�lD.n�fԓ�"�N�q��f�ˈВ�*l�(uzA�/d����k���jtb�|n��@ԉ�Ԅ����:~�G�W)������i�n�@��L�����?���݊Jv�������M_9H���h�c�j.�!ރ?h��6HD�*�?Tx3�G�����c���{1�6'�DTФ��c��fy@dD�}ۨES���&�ϯ:����[ޣ�r���#e%�+���������o7�$wO"�ҕ�w��<_AɆy=��Ԙ􂾤+�H�xÝ��9�L9��(�Fi��i�X
�ދR�~�~��l�c-�'4�*�
L|���Dn�r�m
 ����x�Fo�RT���=��G;�n�t;��T�a�(�'�Н���t�bDV��h�d^�a�A����:H >Z~w�
!������29
�V	q�옹�1c����x���@��bt
Će�=�{��&oR���fYc0-�O�����_~G���ͷ �ɇ=ҦPu�J��I��aP�����Z%N"N$ �;%�(i��t�[b����@�oxݝbY���w����QYH�Ү]�&%
|�u���?gC?�V�]"Bc�;a5�� �C��{��Q�ؐ8r��:ԣöib���P@��^����͹�P�I&���T�{a�S��U7=�t���5�zXU�RĤ�Rr͛��R& J�&)X��N�P����� ��*�ĘZ��n����m�1Z
e��J�\���lR`�K5�z��*�e�_<�[]%d��uhP��@(x(RW�l�Q ���w�������u��{�L>���`T>�V*�ܳ�  ���hCc{�)���/l��O��T+>>�8��v#[5�Ir���<�eJ;��U>�&I������!�jbt�@�+�h%�Β;����M��<x�=�!v���b�����~��" ��z���u!�k�_��mڽvp� c�nYV�`�ґ.�"���&q�^ؐpN3�����"�]�O'�6��s�6�Pf�A��T�k�K�����zÀ�Y�Џ���d��F G�S�%���'P�J�� L�ݹ�c�Ϭ���O[��U�d�\L,��iy
�m���jBX,J8-7<�e�-�B�����Ҁ�5ݱ$�j�#t\{���ĺC6�:����[��]�M]�Xր��Ȥ�7�8� ,P.����}�Ad�^�w;��_���I�w���	�>K ���8���G�{aN�b6�e��~���%�)*F��/~��3"�r�j�"�t;��K�ZŬc���R5蘝�$?��w'̝��S9�����_H��al�x+*/S�#�	����2n�|g��v�C�kʵ�p�l����Fl�r�[8ӻ�r4��vA&�~�Nӻ5_��^=Q�;
:�;�խ�v��1V���V6���r$�� D��CO�7r�OH/t�͐�",��C{Hx�6�#����u�3�rs�k���$���H���	����X����K�2�E��#�(��Iee��;n;r���\E,�I*���=�Jj�hGOQ�Ԗ�2�vƶ�D�2Į��,n� �pH�-��gn��*�xA���~2I����Jh^f-��Hxw{�?M�g��Arv��IQF�)A���⃵��!��FI*ueN8_����IA�r��%�X�	&~4��/��}t�/��� �tr(v���h'��*� �%���=�%MYb�۝� ���1^Y��?@gv �}��t�
�����THo�T�Ա4�d�u�oY��� |��T�6N��u"F{eq��0��vD�ˈb5Ip��胧�~(��&]o ����f-���^}�0w\D{����k�4�������_���Iͅw�ky[�t�? B�$��`2z�\s-ΠO��������iAM.0*��V�30�a|�`l��炍SҖv�<c�������)-�<d�Gk?��1tC�f��+0�%Gi	����UU����$����<�j6��f��hTj�Ć�V"�tݏ��<�y�ˏ e�,�����o�8v�WF֙_�q!�U䌚�0{��\��}�L���Y��]s��K&����������x�X�/ٴy�
3�qwL�+G�P��FE��o#�2NPiD&_�(�N7�c�Ex�~�Ȉ��k}`̘��N��.N��$H�����f��o-I̠�j��N���d�NZ�F�#(y�ܯ��W��2=��zd������4�}?���.v�;���MP7�Op ������9�L�I@�4��"���;7=��D�]�*����EE���0XQ(K<Ϸ5˨�C�	5�&�oa��0.|Dp.'�J��a����C�x}�>p<���gOF�̣Yt���~c`�W����*!����i�0ω�Ά�1����_�-��޹��݆y������=^��t��q
�m�HT:�e��f�D9S{A��ǵXp�F���Qi�Խ�� ��9�c.��<YI߳��Ѡ�� @)��:� �1-�����=v����.�p�)�R�nλ����|!:���ĩ\�}o$��� �U]�ˎ ���z�V^¤
-�J�^/�V ��I�h*J��QT��܌u��6��;����+�f=� L9��C�;/UhM��j�.N/�r%�ɺ�CUP*�Ȅ�;+�40M�K�/.k^y�8%CCئ�S���&&	ȫ3gy0�8Pn��}��Z�?���Q�Ḷ��=�]YN>K�h}C�yS��$j�y��3}Z��|�) ���~� ��ؒ �|��q�9)��H��i�V�9VCg��\9�s��zy8c�c*q�v��J�@5szT:��)�1��ZT� �7ǯ;r��j�qѤh~�.��A��\=�­���e����f���I��(eW��a�+����R�H���9*�S�����K$%%�h�����Λ��ԓ���W�Sq���m������s1C�7/����e)�q��[;�B�R��8�o�۫�Fx�@�߄�#��=����XV2Np�e�;oіDn��m��G���w��Iv�gh5&�#��
�9U���D�ܓd�=<L	�G�a�Й�΁a(�Qʼf9-)+�|�V�6l^|n��%�Q�U�*��:7w�k,r]�%"�9C�����T�� ��(����'��Z&���_uz�����~	��xh���g�'�>
���Z�'���An����}�xk�����y���h���bu6T,"Tڂ����G�=P&�CW	�hM>�lC�lM���4W�3��.�U�tЪ� ȿJ<�i/Զ,Y�{/�%�.*_�w+/��B4�H^pȘ0	� k�(\�NGRD��#��2h��X��Eq�M�o��9&@�k�g�x�O��#&�돖����+&e#���S�Bn�G��ח�Ќ�_�4�8�»� ���p�Z��Ϗ ��шQ�|f����Y�XyVW�^c�Ƴ���R��pv�B�� �7.%R�d�r��1LAhF(��2�U�p@�˳�k�Ֆԝ� ��
ˢ�(��j\䜢~���+�ٵnD}�D����:;@��B��/����]�ц17(�C���}�i��'�Q�r�pD����dK��۝২��E�V~Z�C�W�.�IQg62�}0�6��P��*��iew���"���"�n*�ȗ�:�~��C2B�RX��bu���`eQ�ǟ���k�d ��s�Y��(�tO��9H�����o _
|-A�����H�	%G^�Hm�ي`$iq�(�1vp�i,(�R�5��"��ݲ2 ��	��L������@��1)R����54�Z��g�!>��ٮ�]��ۛ��
��;������E��<)�WJ֘/��b��F��P�[w�v�">"�7Y����B����E�5&�5OPFP��ŵd"���q�Q�?u�1���T�n�K�$�3�)�y�b���r�X��#�.D`�'A�|vɝ��ӵ�$9�a��06K���v҆��bI`5��*��M�I��+A��u� (��t��퉡������x�U wg�=���s6�Lp�8�e�ǌ�����*H�f�6揁R4F��9\��s5�Sb�p,�	�������z>ڮI9~�#��XoV��X�!�k���s�n�B��,���U��dm=}�a%�����������hS�<�98S�S(��\Zyc����V�TA� ��2����w�O�{��Vh8�  �U#n� ���V1Ixzx��(��b�A �_s��d�f��S
�k;ҭ%Er�iώ߫��['����$"F{�;�2Kb%q�o:� �T����z� R@�̢^��Z�鮺����}퇄�5B|�F���P��=��f������minՃ���cNZ�PX�c�N���9-ʱr��׹d���r�"�F��,>�T*��W��U�[j�)�K�S?��|k�ݭ�8�PQ�o���n����?����(Ȧ�J���c�Ѱ�:Vr�TA.��8W�'_��8�f�8+.�Q�f�i([�V�?�lh¾
�=�*54�&A-��2�$�Ʋ���y�� ʜ�
�9��/?�R�oV~:^�iF��bp���-��y4�sw* n]E�H`2p�b�-���������:\�;��[5��!J>��XJ��b#�'��X&�#|�JCjR���[�"B�,;A�=
 ��ބ.��I�L�j)�gg�����/ޏ��-9���v��J�����Bm�����b�=Ӿ.@|2����@�$zy;D�r�	���(48ς#���d��u��=�1�B��7���m�T�Ԩ7{4gT����� Л��A�4�>+MS]{D'}���a���d��.�o�3H��F��[a�v�HL��{Z�����O�jQ����Rú+����e����ܡ��6B<L���;�ޮ �"BD�q%��1������C��q�=ZyQ�Ca�'��$��#�;~h7��1GGMGYE���6}�/��N���t�t3"�wB�#���\KDf�����Ԣ�A%��k�6}dr�c�=��I��Pd�)8+c�Di�Ŧ}���Oo?82h�i�(����B�[]v�
�@���Y�����7@R�L�_ts>[����xA�,���o|7�B��})K�6���D�4���>�T`W���5�eC��je�hg��vZ�2T�ں%�q�	
ll��`Ƒ�ۗ��$�I�_w�k�����"hDH0��0����<΄���֓��B#ߗM"εWvO���̡�a���c�l�;�9hT�`��֫ƌ|�e�0!Q�k"iD� VE���%Á"7� �&���\�C=��qؠ�� (hOW�jꪴ�Y�,mٌ;[w��=���L��=��F?^S޵����B���,�����@#t��)ลm�i��$��ìa����w�:����ɻ�xC�,k6;�>�h�n��<I�Q𰍕E؝<�M�?�|��A��|̶���@އ(�{Z��ț<�88bF�i�zX�������>SE/�����V'�o��eeM�3 ,�K��&-<yE���� �?�ƅpa�cSju=���
��QOg5A�6�A!�p��QA�r�b (D��$��#E�`mD���M#t�@i�L���h8�7>��7HU(��Z+.��w3�ǝ�CH��b4�mF�{�]�*ѯb8�=�b��o�Lp����Ǳ�{�a�:o���K<��[������9�8�ț�*t?|��rc��6��
��B�(۟~.�&�h�d���[���񭥬K�_!�%h�M4��>����������ŏ��`u�6%8I�7�(���>�7O�bv� N�j�xb��ϷA������KA�Iܣ��-g* �O%�m�ͯ�H-��x[@^���$���R������t��'�=4PGx���8�Z� �g]g�11��'L��=Y����q��m�4�q-�T�<q�w'�m��~^Pη��_��c6��Uqƞ}u�T�� IA�R�Got��|9�Wmx;��o���'~���38.��ǻ/#��f�8�Y�b��z9Ǘ�H��l�O9���z���"(�e��┴׍O~/�U5��^�NY`i~&9m�1FP����'�1w�S�k�|J�S�P���Pai:jk�6�y���U��7��D�2�Y}P�=+D�]k\�S� 5�ˎ�����t�%O*�GQFj����7����ed=�����r5�[��Q.o>���c!���믺��D6�i�!�����`��I�	��K��}��-��D:����$N�L� t&��������.�9'����['��ُ�w��LZ��={ֹ%')Ż>j#ĕ��~��DP��.@6c��i9i��#��\�l!����e�]PыX9�p��v��P^M��j&����G�f6̀Ӌ��7�2����o��ﯦ_��5x(.4����D�>}�Ȼ�|O��ܫ4��nKR���D��+�#d蛆�~�X��@m���AIQ�
p�&���ѓ����#�~�Dw!k�[x�P�����w54�Xܱ�1c�v[_��v��(R�����A�D�&�!!��	4x���]����lr��w��s�{wX�	>�a1���e����������S|_\S�9GWy�>�?�p� ��ݹ�Ӄ�.�(��U�ď>9����ُu�b�A�y�k&�;�K�Z���l�O�Č�k�8G&/~��~Msxy �'�'M}*�a��\� ����"^Y�i�}�R����[q��b�E�P\Jt����j�#����@v��D�q^-�	��7��\B'YxOR���$������w�X�D!�"�4�)��a=������� �uڍ3ڬ����Z��r�v������������=�s?���H�,�L��W7X2���|�r���X�D	S��
��c$�v�ƞ�--Y�z)Ǣ7�� i$��P��	+|��X-�:��LL�Z�U��X+�M���'"��U		�w+���R;[$�j+�-�F������:��#�%��f���ܞ�'p_��>�����q��|�z��B�Us���$Uy��W�i�-�r�Y�����e�٧�9����V��B
�]^s$P}�C9�<̘_ޔ��iA��ڧCx�>�	�����g+�pUN�\R�����3��Ԃ�f�<�k�|��R���PM�)��M=��
�lN���e���Bn(W�l�4q?T�)S�2�${��A?O������m���tV[�KDš��eО���-�(Ӓ�*f��ԫ��t��6d��ۧ}�~u�
��D�ˮ~��b���I�"^�-׋�,�E�4t���I2��|1�6|�QZ���Z݅׿���2X��&�a�02�_ I������=Ez���D��F2��wc� ,�*��fQkT2҃�"IG�� �X�4N�5�&��	�
�Vz#AZTr�_fz�����-7�E���3'V��;��H0��,au7�l�QM}�PzHY�!�	�����^�[Y��Qk����K(Z�|�:��x��Ow�x��w$lS�A���׎l���W�h�����m8�#�33�E.ҌWgǃ��Mw�1ӾNV�flի���'a)�����ϱA@z��q�����o���4�$��1�鏨�wd��'�?z0�V�:$�,�X
�!��x�\f�=��S�l�؊!z%��4����`�!-<7�;l;T؈��>�E�	8	!&Np�g�=
��rp�=�f�~��$WE� ����2��Z7+Ɵ���%��p�\����]��n�O i|�݄�����Y��} 7��5���W�[��D�����c�T�"���¼�*T��R��[ ��]��L�h��~,�DO�Z���~>xP�VE9�dOE�a�� S`�2�oL�0�/淸���$5������O��1.t3`Z��j6
����4��iJȈ�OVy�P�\ڴ�Kr�P0D5e'^V��+ ��,e�5��T�[ ��Hfm�٩��IO�$>��S������Sc}&�x�ڶ LJ�@���E��nG�bDK���ZfНT����g���zsδ��I쎭#m#�4 jr���.k���2͒�]�A�L����oぬ�I�0�yMV}۳�q�P�����.`���a,F�!�H��M�R���%\�&��O���M��)k��Q�a|J�y�۪fq������e��I���m���~�\��W�vSb~��3�~�5���UY�#��p�x�KZm�Huy=00	�E��>z��sB��.�NGe��'?��;"8²�[Gm`��L2Q]H��#���rx���}&���z���o�����yRow����lcș�k��y v<������p��f�nc Do�>��[���mCl52�j���M|����5i����<�R:�}�V���i��1�ÉBh<r��Eq����� W
�t��'c�I#�7;���>b׺��	�/�|[�A,[�����Q��@�M���X�L�r��_���6:(L�b�����q�
�=���� tIF�F�G�]����mʿ��4����~����n�2��U+���~�)%B[ �Na��L��$�\��4�?(��O�e�b�}���u�-A������f	�0�R����m��!<|�?VD�9Ď��P:�S>a*�%A��{�F�k.Q٢��wj	'�q�:���󤯚��z)�\}�3	�xU�A��c��]8M��Qj�p�����ׯ�@�Ak�9 ���Z�W{Ʌ]؈��� �)��6���_)6�`�-[����Z��ׁ�~g���쫃��3� ��B�wO~2Z���)��H��m�N�Oz�))0"�������Y��I�V�n��P�:�R�
�$дِ��/��i%_l��c��?����K��H+�t\[��
�fz���X>�4$�*���hG�x�7����ɐOY�� �f4�aG=�U
ψ87��D�]:��\,����)S"��\��s!�X}IY^׻格��&t���IG���8��b����ېsĦ�R�M�z��OzFGX��ܿ����,A[�'�`�+y��q�ۗ��Fu�0�W��)����6=31����|��N�8������۔�b��Z�y5�"5^�q���b��
�a����k@i�e�1�㮢�3/�؉�B�_�zͨԶ��^3̔|�&K���@����7�߿7��`��M�7��Z�.�w!s��A��%��f��U׬ɻ�
^�<_P4����.�z�a?^aU!�ο�Đ�a�	A��� ��D�	|eB���Sέ<�:�?);u�'�Q�O����r]�D�LykW�f�%���3�� 7�5?��0W�}܉5�pM��ұPA��������0d\Y�3���$�����~����4�^���r�jN���:�o���s�8�L�'��)��A>�|��9G�����5�Q��)��� �<�V-t��>Fx � a�'Mǥ�*28��vxxQZC�Qt�$� ;�X%ft#�a�=|x!�!n�U�Hg�d�Z��Xd�6�E���F�B|
�oɰH�i��OT&2$nHq�`d��Ӻ<��G Ĭ�\ʏo�LM�D(k�f��c����ax|�\b��y��x�J�6��;Jfht��q�����z���7�M6�wVs@A�l��b9S��Q�V熻9R#>�?����S�o�)��V��j/�|�$��̘҅�l_�R�`�ԭ!�DF��"�4�W�0ۺ� N�hb鿮���<O�R�̤�X:a�
P��d�B:��1��Vc���u����)�?�h�8�?^`5Ì`l�+�|)���?��WQ*�L��ZRf�~z���O'�����ep
J�*7�Z�dg�R�����<Y-c;@�3Ռ^���I�W��%cj�hYJ��)��JH��C˺C�ȩ&j۫����/؋"��H�F.���%�<9}	
l������Gp���C��x]u�!k�s��YM����#H�tm��\W'ں_ɹ�g�nV����ki?o5;z�̌�aD[y��
(0R�����=}�>��n�a�\�K�<*�o@j���=7Bx�+�9 �a��KF2�쁊�oI� �h.�%b�'~��Ο�`� X�9"�W2s�|�� ��+Tؔ��m-\���>V8�����]"$�p1���>W��oGj6g�++c;�c�F�qs�ߩį`}ȿ�:e5�n�5E���p~q'�������������ay�O��o��sxY)%�<�ނ?Tҗ�`T%�� �?�$\�O�p�Ѥ:=鬕YXB`_U���^���']���<��Y3I�G&>_9	C(�̫��gr�Do*Gz+BtYӿ�!S).���Y������dg�eo�f���e��bd<�q�(��n�qqHX��)�T�A��	i�{93/\����]\'�����AR6���?�6�}�+�:ԗٔ�?��O�%��D��Ug(%<N��AK�]�_�啞��
eKs�*Ks��	��p�$��\fVt��!'kz+����2	��^bU��2
�7�Oi��6 5��������<��v���{UQ�9C4� Dj�R[{�&�ܺ��`��_]��D��'�9q��O���te] �/��'Z�ᷦ"~�A���6*�P��&F��z���W`c��r��=��;��ެ��8��}F�G	���+�,�'�	Kr���0ɿ3�����ao��DDq�ʣ��-2�?�1��E%@Pd�J�\��Tǫn�ܾ�9~9lYʹ�g̲y�����A�����_�#Wis��4��(Q2:R%A�3N=�B�_%L��	2���w���#�#"�F2���f�>Er�����G�8u���v��!$�T=nc���v$��j����I����r�i�?��S�Q{by���>��E�HJZ>�`1tLD��!E�og��5h}b[L�.)H�;�̾S�-�L���|ː[s�b��z��'[�J�	��~�n�؊��#��x��"����<�t�?TIS��ߛMh��8��_��Y6�B~��9	�c]�I�|e��ǁ�:��bd�
�>�� �?��6�4d��b3�s���\���Y���{gf�����&�]{럻��( ��l����/��I����7�H�#��Ge��?����i��u����*�q�k6|��`L}����$�Ή�+D�8 ˍR������������; ��U�~��9*� ^�)�[	��:OuChg�i�vx�)N��Y$�� G�F"���TE�P���UyI�������Z�6�8�ft�%AF��N~(���L�q��j��(e���^���Q�����#�o�Ʉ�ҡJ�iۮv0�m��^��Zw�w�`۠/JX�����!�(��:}u7נ�>��r��&
��G�h� �h��1"��h�<v���F�-_㱏�	���:c�v/J}f,糩+ҵ�4��};4�)�~^�VN����۠ٗ�����T���n�S��]�\њ�߬�����K�j�`f�Z][�H+�D����9��D��T`�*��	����|��%�s���^�l?��D8�������(2�/�bP{y��t�K��Aϑh��a��4��O�5�v�E���Y4������{g��	�U����(�Z�Ӑ�G�Zc+�����̃ަDR͒	UL�N��"��%v�&=��݁{��	`\���+�C['���L�s{�mEf�. �P�����n*�b�=
�� ��� ��Z�[�X�iE�Q$?xHÁ��m�� CR%��*���I�5\/�kI���g;�*D��ԁ8yIC�
@��d;��A���*�\�!~w��g�|�1��\��6����nj�ŗ���}mN{��;�B�8�1�V�/e*�q �}	�lX�_���*K�E9�;� �̥-�x�[=�zl�Tg���BLE
�	��4�M�Lplk�K)��ʬ��x>�
^.���Ld9ЌL��!�3P��@=�� xH��%�*�7��~}_٨�;[�v=ao���� ����"��=oQ/:�ݶ�����?I�Gy>I4]��n���k��ñ�\��������2^dK_�j�5._�q�at�}*�-���Ÿ�*Mbɨ+~�(�̈�W̾�BE!܏��J�\��v�N���G�?wwCdv[N�{�8��z�W�\��cga9�(K�gQ.��O^֡��\�Jl�Q�LY��G�y��$w�gbܾ�����]8�@������%'�����!^t����[�?��4%@ع$
b�y(J�0�& *���Ss�ԍ�8<0�}3��9�ĥ	���OY��x�N��}^�s\��	�':�n��i���Xٱ}h�����jL�:���$ Ԇ"Ў��f���\]����g	0�p��e^ltx��������I�4��<=���{^2����	�Q�}�!K�'�ug}-VR����dہ���Ͻ�q2+�#���t���.��k{&K�}u����������y�5q��:D�|"��aO������=I��0$A'��VʡGx5���x�%��`e�ް��;%�#dl�@��%�Xd����yf���<s���$����F���K�&%���wyV,.ݱBO����0��3j@~e��N��D���WK�σc����!Z��{ws?Pc�j�G�#l}�(�,�f���aI-�"�����pU�MX䎒�xǺ� 1y�ɧ9�w&{�$X[@�-0ڥ�/Ax��\��׋��Q��"��6RC�}� ߻i��Z_� g,*d�����;���,6`pE~�����$�Ю��Yc%��������|O3u��wȅ�XB:tѯX�)S�����0g���s�3g�3k^�"�B���65Ƶ�`��%�=����z(�ء!��V��~I��P�jR%���*3\|���7꣗߲����v��8w�ΆD��?Yu�)ւ�r]��)f�Yq���-ѭ��Mz�/�`k���s!��1�˓Q.���z�
L:P���A*,F�Z�6��ׄ;\3��^!G�����z��7d�Q_.;՜R$�%׉�m�������/�,�>�\Ŗ���C��{v�WtbNvD���7�{)�������Œ�5��/���6y0R��00/�Z�{��b�A�ʾ ~��#7ELFO br����$`F�?Y>�U�s�3ϻ]E�
kx.�w*FP�pT|!G��.��q�`6k�P�㏑���+����������ml�h�c^�T�qZ�"`u��X�Ss|�e�k�_@H����x=��s���X�kK0�Y		gH{�J�"��3)	�bFJ��[IR����P�a�*���,8%�]tp�ڷXp�Y��O����2$�w:"e��+l>���[.e�P�+~��V�{m�:��H}�-w�!1�0Sv��f�� Ѓ��[��|���*팏_�)���º	t&��P�j�7��@)Ð�h .���r<Z�@I�L�;�,�/÷��d�l�81�`��ȧ&��(��a��1�^/%����;.�+��8�(����|��]�ֱI��	��cݠ[-E�<��
U��C�9L�Kgy��Ԟ�3�@���������\
C��t��8�ƕg+l�%�Fv����$����g�|��*�-�L�\0(U�9����ټل�c�Ӻ����i�)����7���'t\Ѵ?db�Ow�:VJ��U�"�y答�a�c���0KH9�-cȤ��:K�8$�Z�5�-�E�������G�令+fj�x`(L��#�u�_��⌀�!/�d������\�Xz��w�T� ���/Xu���{�v��b5�wcN�	=�]`)�uer9��\��8��f&n���xT�-s.>�Y��?!�G��ǭ���4|�����F��9�� �J*�I�F�pP<���;�IOd��4+�'�yM����$f}��x�'�t�m�=0Je7�?tk�_~3�y��bzY�.I����c�$>����������S�*�pԾ��/�3��F^j\��g����>�������<�pdlgE��s2��Rb���m�ȫ\��B`|�#=6a�����E4�3%���յ�^BҰ�D��
+�]�.�Sk\����M�t�:{t�Z5��F�%_�a��Qi���C6WV��P��#&�W[jc���%�f����>l���e�P���1����?�E�)��ۧ ٦��1�v��М~�j�Pe����4��������R�j7�:B�lt�-ƌ�	|�:*w�8|���}����94��].!O{�zЌ��с�*4n��\�kag�Z�;:in�cB�\'_�!m�"E��w�n%ۃ�uw+A5��=�{4��s^�u��6�؏��'�����j�e��'%�;k��E|4K$��!;yDh'��r+ĮJ���棔�λ� Mgm	w�i�(:@�"[oX`<����/[̒^ǫ9�y�ao�L��M�?[�;!��	#؝0""Oh�3z:;���c��a& &V*Zs����ir�V��6i�S�t%�;�1L�"'���Rd�FcHO�"��2&ZxLDL�ğ�5.���ޅ{��ʍ�<`��4xk����9�ו�W��)V�3�Y�5��/��jw�lۂ�a�X�a��,	�l�K�rSJ��Ң�"ay����6�H�/�ʱ�O�~F�P]�u��lݓB�+�ʈYש��U*}T��]dd���<�����}�lm�$H����3�d�����~h��u��ٓE�W���)b�"$8��<\"���XQ@�YA�!�ʀ�P��W�y���^����N~1cC��YP��P]ÒĤ��2)���Ӟq(f���3���!�j�;5�����&4>T˩R��`��ӐC���#p�]���,H��1b& �_���v�t�<��V��و6��B-�m�&9�gj:������\��n|�r��k�)�M�{e3]�='ᐓ&����@$�ǲ U#WY��L��Q��+�~� iQ*��sH1��G�E*�R��1TE�޽e�E��Ʉ�"�7g�t���ݚ��˥9��ʜ"���) h}��(�y���5�0�W�d�t�w��Oc@�(�د6�3mzub�Ӵ`�ϑ�	>�lܸ"�.0����U��`k���5׀����� .ej�t����; $-[G���6��>���P�2(��ϻ�Q"4���y����d�#GX�(l� b\������WSV���ߕQ�b�cjLy�)�M����v��]���'?�	�̻�$Q!e�2l^E��"OGn*��i�
IL�f@��ɍ]���Ӽc���#�1*D#��=D���	�u�&z������+t{�I[w
4��(˭����1*� �a&���x5�3]���5S�,�yε�l��M�o(�D�nভө֓��/,KKU�陟y�8���E
K��t���`�*�e8�Y�t��Ԯ<3���'��j,��ll%��s
U�3B��i8Q�J�
lೳ޿sNr�(��h�cp��եU���E|n�9�(���J�{�F���d��/!{��;��b^��У�w�y���c�}��d�d���XؑA�
1 uq�8��u�>2�iNÌ�$T�EZ�o��,j�(3�0���K�
�ţ2�/O��h��ƒU����7����G?~�ojlw��Ū��hVNH�B��y����KP�q7�;���J�[�i'gcVm�͉Q�͙�����Nu��Y�1�r��U��҂DWyے�
���S��}�?�k���3,�- ==^Ea��:��'������z|l����ZīH�M�y�^��B�*�(�ԑ}��:Ü 9��	82�e��9�.P�t�'�.ʰy(@�+�}Z�'eh)�&iC�8�nEi�{���W�*�.D�?9R�Ǡ���Pa2�H���Q��:�8n�� HW7��~�$�N�Ƃ�2����:�u�V{�y*a�#�N��R�VH�3���$��#i_dPn�*��s��u���.&~}��2�<�eɶx�k�6Β<V_xQ�/���/O#�@���'o�͞�o���D��+e���`�t	%'�j����~*��q�Zl�40��� ��j��]��B4��v@:�)�qXK<�eF����ևZ8t`���	~2�e��G[�.]p�h)$ܪ{93G�`��pS�����g�K�(.0��ٶ�A$��sF��$e� �+ ��q���ưo֫IW5-�X�4�ƻ��28-��0 b����-9�e(/�x]2��އ���|@�.B;�Vd��
�*���9mX��\��������##H���[7��Y�׊��O�.���9͠����t����q!v4�<��p�ȩLߊ� ު�*�ϝ���ĵ9K]L�Ͼ�v�aUF#ݛ/[E�-�U�85c�'�̧�! X�omNJ3��q{�;/���V�l���nK�Mj��ḛ��K�[�鴂�5�J,�L	_{~U�]ڱ��9]4ۉ[Xfoa�έNuu�V��ʧ�dl�A�e�����A�aRd���Q�;���]/`6�mc�/?,�W3�3J�f�?����15��� /�K���[Z�ND�����YC��9h���������9�ݻW���łE��ڊ؀:����d��� ��/��wQU*\���K)XWX�F��4��H�SR����n�O��YΞ��%^}H>�$����vT��=�f�?6bK(���Yc�ѽB�>�^Ӂڼw��.d���A�,�S��,��] ��F_C�+p�Uk�"�c̼������Q�~�P�x�����7P��U�Q��Go��2f2�C%���wo#�Yey�K�Tn�F��"p�y�#���S���c`��g�4D�*S���{��Ag�2n��i��>V7�|�{�#�χ?\;o����4�j�c�h�~�f`���@�e���)�H�ޑw��^��������Q���V.p�݄B1�Oe��_�\��j�3���׋�hĚ���9,�;mz2W�*�V���tN����S��v���p|�[��~*�k�Ja�JJ:J�>Q�ARC	߮�v�nAKGJQ�X�1�3��"���B9��ДU�%���m�O��:���T�$��2N�D��xE��+*�=k�7q��zN��,r��}��GB;������D�|�7rv��mUO�u&"���J�C��?(���~>�Ql$7c[H�r��n\�|��Dbڟ� g��z���|בM�.�sG'�������_%���K�VY����z��)<p{`oL+͠H�Y�#���v�%��Í};�1t=j�<l�
�M\P6�4܏��}r���X�l�f�d~{�8������B�_j�ɢ,��xF��uf����c�Ƹ�U*۹4˱O���
�:=�'�
e����o�d�=�e�+vܖ���,�nI4w��u͛9Aɶ�]pշP���%m�̕j6u
�u�bܑ:������.��w��(,C����������%�)��3�)�,�&�ptQek�9f��/���pdK�j�c�8&�85 :e-`[�����G�[���z�$,�~�پ�X�g������*΀��7�p��o3ݳ�nα�z�۸��М�s���*����G��)�qU�&D]�������8��u2�i!�5W��jgQ{��4T����Խ�I�Dx����=jÍ&�[��~d��u�`����s�m�����[@�Ѐ��4�0}B�9���Y�	�a���"�����|���x\�cO�X�h�4������{��w��x�ca�.������P���1�e�dF�	���z�ܤ���j9得.�������i����bHz}��r�l6��L��������6Sj��.��Y�6�c�;@���E�7���N;���	�UFDR��e�s�F�h&�e"��~6r�_�'2���JB|���e�q�=�08_ۢ���o[�8��-)��BU����ǐ���ۜ
w���2M���Q wdhqS>���3)�e���ݽ�aQnG ��Е̣�b��je<�-�xB�e;�V4n��6�X�[�	�s�y����-�,T������8�7��JgR�HUdDH�zգ��H�i'��O�I =��Ps���|r6�U�Fn�a5�T�A]���!F�E�h0��X@r��H2Ĵ*+@!YFA
��'��<�NO�TӨW�*����(��}"��@H�W*u�v�*���iQ�аg�R>�U��v����W�J۝;�J厯^}�`������鸨�r��D�|��4�Μl�i�_o���u
4�s�=�qas� ��K�'��3@s����M�����a��*��I^@ �A�y|�ƙ�.MJ�W�}]G���r"�1��W��R������J��w��ŹZ`4�|�Zu��,���B�A�u�"��R�3g�o̧�N�|Zy�)�[i��Q`�J�ь������h�*T(��|J��ȈG��K*?v?�l&�������
q�}�Sl;d�ׇ~
��;�Z�:��,TÉ�q�$�y�f/ U�.ɬCٍ��[k��v����H r1�RpD�%o�vS
���~���x���*�����[ԋM�^�#�a�-ҺO�b܉D ��nop�\���
^�8JLD�c��#3Ƅ�W�u��s��m'�~W%�� Х�
�g��B\t���JJCa>��łO|��7A����K�S���,5�!���݇(dq���nn�N�f7�:���v`k��6v�99�R_>\���ܘ�MD�����mj�k�&�YںMY��o���[Nw��6Xx��~��
�2�C�MN�;͡w�<�zJC_Blr$�Z��>�W�S�^kɀ�"���k(�
�6leu�%�f�2U^��a�OI�F�e��8k�h�j��꺻!����bz`Tˬ㣙��b���&��ƭ�.���oX[�ij~&S����Z���������o�n}�����B����G�a�]?�X���M�ˌ�·�8HI�+mBi)�N�y�wBk�����T��O����Z�p���ς���m H�9�|��ok�	s릅����l�ir}�a�	��f�Si*�kZT�A��O\�ț���
����[@��jp\�)~�,F�H�H����#J>	�~G=��䆠�J�<���S�W�U��w�sa�u�F���{�zy�h+�`9[
N� �3 ȊW*�؍H]WP?�&��`�w��AK�;���
��kV����Ξ�D�n3O��k]�Q������<v����_]�yjS���,���'[ȟ'�	ZT��x�=m�,�����sx�m$C;ƀ����C�������@�;t����1��
�m�B>���a���P��(�V�@x�-e���/�j 	��A	����o���X(�R|r���W�V|�lfϮ�޴��d��h,kk�9 ����GE�CkWZ"m6dɛ��Po���o~d�Xw���<�38R���c��2#.9G?�u�}����p��I,;Fp�#rqT�%�e�'��`+'�I6��MG`V��] }`0��UG� �y�{9�<"�i��|Z&Ç�ɏ�T�[*Fr/�"a�.CM���O�/�rT�=��I����6f`��␾��p�O5�����}�/���N��+�-I r[�CiR���[XR��V�~�E0 XDw����JL�\9�:4�'s��>�f?j���<ס�_[%c�
i�0���-��'��4m~���A�B4�̗3 +�s���[�r]t�0,M!�Â8�ʾN-��v�V�+�g!���ic,T�k�m�����S��Rn���d�#4IH��W6�wTJ̀<�ϐ���a��u�It��u�X�=Q�s�)z��W.&S��@.�o�E�_��]M垁���J�����)�b�����tK���%ív���ƭ,�p ��^�!���p�.ή4$<dF\��L�fe_�y��O%; �)w3Ǹ�â[�QY�w�#��x��G�%�����?�UŃ#����L��X=����	zP�To��/��h`��D��-hC�sG��q�(a"�#�� A�2��C���P])��V����҄3�+k�쳍�J�<輔?I�xO��e����Nh��!�]h�a*uk�k<�A���ѷ��/ha���d�kh���~��T7'��J�P�~yD/}�2���1��h*ۘRj�@�Q���y�3J��\u|ɥ��L�q^[�OG�\��P�vD�ME����0v~e���w���.�(�����ogA�=�Y�*�c�M�:�Ē�)v����C�Z�$]��1�ȧ)�T���67�E!*;b��WO+���d�9*��t��(�LH�s�We���A�nM�qv�EDv���Pz��e��C�DA ]h��PQ��62h@���G�n+�m���;�[�
��m�����
ߚ�A��Y�ā�͊=<0m����5�Jc���J�̂X�g#��9S���H�Ye�o�Kb� E0�N��(]wJ@�s�qE��>�6F-��_~䁩����Fj.�k5rY� �����H�C=�o�P���:��͐�wU��sЪ������ʼ5����"*0�����d��ն�@����27/iֹ��vW��� +��{HmM�� 9{��o)7Q�[�
M�G��s�uLe �#p��)}�a�Q� ����E�E�[:�`H�%���Q��U�dR��ځ�c��Mn�|���� ��E�Ba	r�y�<v[�J��?���@�r*�I�J$�"CrMo�R/h�9����t�?I��P�S� ��xy�Cl�T��|DE�)�������cQ��f*��(���
6�Vbfz4��Qw\��kH2t_B�TKX�`�[۱���C�a�.:����U�<_�`rE��wD��Fڐ��jT���|��
�=��6�ŋ���;b(0'�LLY6�Tܵ �^F��Ѥ-���U��~}��)/4+�g/?{ ��@QU
���)qftQι���+8�(�[����<3��~j4��I��:M�I��f�X�K����QR8PHGBdE9'�EB5%�HY$��pr��XgЖ6��C��]Af���<m3$�V�����>��+2��&Cj���fǨ�`����� \��vf �N5�q�׺LQ��^T�� �!mІ��ȷ"�����/���,���1�:z��<���E0^Xtё����L6P%H �';u�����j�!ѩ��G�������c��}�3�%���X]��b8ko�`p�=�m^¸���]<��%�A��	���B]l�i��G�4$I�Iɖ�`k��������Z�*�=���/6��ѕJg��#�Xچ����5w��Ų���M� a��H��e?�91�<�Zg�[	JI��m�Jኲ<ƷA��+@~IjQ���u,�!��u,-i���^zw(s'�r-�]�%������S��hdHn>��Yq�':�|eNڸ�[��k�}w��Z���N�F\��;���n�'$�P�������Q�:l�Qn�Xg~4��i�/��ɷ8��z�FY��ZUI���!0�������x���T��U��a�$���@�)g�ЙS��C�.[�c�vk��a��VI�&���T$�:�n��97KQ��� ��7�<��^i��� b<S�ȂN��M�d�	������?�M�w&�ۣ�B,?�8x?�;����[}�l����u]/�B7�bw�cx��u٤/ك��QuNJ�.*�|��&�.������w��æ���Z�)�+��K[Ȕ�غ�eQ���m�8*�F͊����~���ím,��St� Qq����
��g�-�� �%�Y:��%sj�@j;�&b��(h8�(T�_O��c�(fVl���^�or��<=�3���Ȼ�����+�Y7�D�d9;}ZK���0���zm_��"P�q�>��{�Hq���g]\[P��Cz��7-!�C�����G��nT]RW�\��� �eJdS�1������~t��x�5Ic�iy��� \����*��y�϶F�{�2� �^'P��y�i:��v#���n�{��|���%MȦHH$��g��j���1���V
{�����ܼо�im���W���� �V�L:H�����B�{��M�wk7d�7G����;��]L�݉��e6��V�]���J�;�ՇO�������Г�*�]'>H����N�l��獥����7�����U��\ڞ`b2��Eg��&���m���
���a	F�:֜"l�����>+O�Q��o�����c��\�j��J�}��h�?�:�|��@�k3�<�G �].#�1�}&<z7��K��ɜ���HG��S ܨ���.�*V�6�Uo�N8V��9,t�m[�Ge�ʈ�֟a������P�}�3i1�>j��hcE��Zs�B:S��TD:{�΢6�s��������}�zĩ��*���#�	����g������	�c�	��+?Mcrcn����<K��|�ͺǽ��<,D1����qN,N�%.��F+McF�0�-N���H�@���|�[3(x��H+���I�,��j'��	�(�e�����@ί��U�ԡ��������g\�l|"C�5����Q]��,>�қ"��\��&zh<,nH�����.�	��R�k��f�Z�9��w����x ���/��8�e�s
���=��ѳ�#;�^<��\����ޢwBB�묨�i�����jq�+j�V���=� ɹ8�뜯 @-�Y�h�]�3	�J3~��χ��H|7!���z����X��yLk�#&�u��_��T.�Wخ,V���**��1Am�@d�,�F����iĩ�'f���y�/D�����@|��	�U��_�W��:��#	lӠ`�m����mZ�;�?�o���J���5y*�s�u
�d%��:�d@i��gQ{�}�_Ċ���U,<c��G`��G�\�����N��K�N�����Ԙ*6���/RQ�g�{�=jО�=�=+�{�E�^_,dQV����W�tt�b"�c䄓�7�D���ʎ7�ۯR�G���è�Ǖ	��/Fj$�Bz�i��؀NՉ��t�VWH���Șe��>�q�g�[�<%��K�ek"n�jV9S\��#�ڻ�$~d��8&�%,�ޜX��	�Օ�de�f$f�|�d�"��.*kX��?��ˠ���� %Ѝ��j��>���#I1���B��F�|���B�N*�,��E� ^Ϸ����{(UsA-6#0IhVh��Mu&=���B'=���ː�>�u���8�����~���'�Κ�� ��J�G.��(�FVT�&ҵ����9�$o$�i�V�{��ߐ�`V�D&�d��C|KL����� ��a�$���[�5�03���ˀ+�h,�.�N|����+W�f�_>�G~i,����<|^��]z'K�{�k��5P�	��
��ˤ`��!�r�@��aU�]��[Z~a��6[>�\���z|� �T�Vu��̸̢v�_38���U�ju��3!z���^��̒~���/����;�؍��+� �z7gBD���'�E��ً���]�`�<ŉ*	�)P�A�$��0�G�b]�4D��b��+'C���SRp�׀�f3:A� W�TA�sOL��]��+��|�h�q{9_�8t#��O5*��ҧ�����"a;�����&(�P�D��}tĵa���;s��0}R{��D��[n�qKIk��c�@5	>@t	���%�5z3�ըB�n��*?z�ͩ��K���6U�L�7m�u�sAc�a�o<zEn�,�U���M�û���J�̢����Qk��G����_%���d���/�FG����WU(���5�9���ըb8Odv���2��VbJy׈
>�&��B!6�h߯��4��?���	WO�m�ki��潨/��0к��z�1�Po�P��s���D�?l�	�]�-x��M�fq��L��M��l[��hv�G�skw��+����;����>���;q�Z�j-��kW�R��(YOa���uq:u�~�?pk�7&f���K'n���D[8.?�O��`HXB{/���_��{J�/�˝y8���#�9_.`�0}C�'�}�~Bb#V�w�}�С����;N�	so�������)��N��]�ز�^�z�O(G ��9
��)n��S�sǨn�E�^�0���v4��Ⱥ�2�L�U���(������Tw5X�}Phjzb�������'yI��f z!6m`�`vQ�B�*O�o+~��(߰t�L68=����-T�+P�ګu�V�mu^p��f�F��}�$Xz�w-sj�p
'�iP���l,�. x�4��tO+I�S��h)V��O͉y����/��,`�+�u��8xi;m���|�,�L���8Q� W�%�j+F#E����>�������� @�XĈ{a�w_39����-�Zz�c��^}�T�	l;���E�zE,�f���Ʉ�S)��E �HoL�L$����_���[
GP=���:u�ޛ'�D��)s�4�6I<����Ӱ��T-��@�:�h�� ��m�X�i4ӣ˦8��s�S�����1�Kf��W���G�ΰcW����޽�t?�EԾz���T���'*�W���,^-�h5�m�m��8|����ơ�������P�	Z_#'���v�UW!��ejt�-+r��wQ��4�1�7�^=�:f��7��m���uh�$W��k�m��U�2�U������>s������]�Y��ї�~#�z�ɧ�H,�h�l`s�ϣ�QOa����s��ץ��N�F�(�Q.�����Aē�pɘ��re��ӌ]��]I���L�BQ�u&��ӥ
�+ʭuzE0����w�>�Eݛ����TJ)�[�w� 4��J/ $�k��s���cWyN�������6|8ߗT(��D?�ƀJV�������s⣍��,+�w�ŗ�k���^0# )��ExHt��O>�w����#� S�z��	�l�a�7�fE���+Ѽs�V��d�{���R\�?�*�2MlVSQ�� [8���k'�b�as����y6�H��X��_�X������P��%AI��`w��!�F�p\��m���E\�5�};�-`Ϛ��a�E��2�6�2|=[�;Xh*lU����o��^���u�t�VO�>���r�+���c�{\ؗ3����r�qq�ZagB�-�gX���|�h>�<̶OL����N�E����eC�����?�/{����m&��z��#qD�z_e�?����P�@lA���*H�Q8��L� �-��Kv���}j����P�5���Pr^K��`�u���iI�%߂{�۲�GD/,76� '(����nt�/�˥in�u
yt���
4�ƃ�C/�ɫ]֤�J���'��W��j�ܖ�V�힄���;��w�	�(;ADÌ4g�:���ouېLG�����=4;:�$�_fI�HqS�	��n��%���&FՄ�#���CK\��zy�%[ՙ
3T�jm����UX��fk>=��2�H�Ƨ�3󵅢����7���A�,Ks����=i=��vG?�j+���imЋ�%�:ʲk�>�ri�h����� �ʨ�@'\e��C2shA��,�Q̪X<�gRسRN����d�+U)o��@�1���(/u/���a��f�Ez���f�7��ۺ=9�U��E�h�u��.��=c�HQ���"旙���0�7b4
:J���_C�����S0�uuz&�s!Ú�d�䵻��,��2�p �q'j	@��OM�(��|Z�/�@@J���� `�@�["p[x��O�YKs���Sͽ�p�%]E���{M��Qo��D؆�%g��$W.j��_�c�� i�u�9�P���[D�m�L����I'�����`�A�>n@a媅bPn
�Q��T1�O�YeI^Jo%����vY!���(��S�l�f7�zAd�� ��E!��\0%ms� -"Q�jH��B�a�keX�ΑZ�M+���X��\��Θ��G����I�9�we� �H��Fv���Cw���$��N��28<8�-/bA�ЦK�C�*s1W�����K(��t#��$>]�g��P�L��5LEq�푴C�jͲ)Y/��RC��M<��5����e���	۴��������A�g�6�\���G���	jo2��Һ4�Md�w�I�MJ� [�����!��{(��?������`gej�"gxr-��e��.�ݫ���=f�)�I'�O6�B�
qI���YmCbr��zL��悀P���1H�K'z��<���o���fQҪ�&�'"�1&�Ը���)�LDA+ �e�#�1�$B�rhq:鍧r�5��h|FpE�<j�%��RYS|���\*��d��_'A�sc�)�
Ê��*�i%$�IVLb^����|U�]�5y�e�\�{��?�v�)�����2O�~��р�GK�:n�|��/%��B�T��7Q�2}vEƈ�\%�Vb.=JZ�yE%%�H�}i�x����8�j�۹p���va����Qp\a��Wd�lz�Q�!I(��wP!�bX4��;m�<^)��I��p40W�O��A^=$��L��or����o4@-6]��4!�!nTX�Y}�m����i�8U���Ж�Ff��X��њ�F�9a�]�pr�����N�f�HC��H�R�Z:�,�o��� 5 o�g�Ȓ���u_-K �W���C>��{����`�����ǿ��{�-�R�Ϯ������hQ|^�h���n�y�HŦ�Զ�6+ ̹�=,��8��Nw%;�֧(Yfߗ2?p������^��-Z��BL�"oע%���͔ͦ�!*�;Պ5��>�g�F,�y�ڜ��f��P���nw�o�@e<��t�������W�4w;/�S�Ǩr��w
�w3�6�^!i>!z��s�,�ׯ����Q�Ϲ?h�ٖF="�t<@� ��,��/�,:�jrM�-5i&���h�� �=��/��w��3��.�
��f�փ	5��H�L�D�s���m�;4I-�n���d��b�l߾��1	�h�%T�EQ��T|��[T�ۛK*\��S�:��=���n��">d�}7�u���d�z�u̾��~c���~��Kelg]����%D\ u�U!>3�0u�:�(���N#" ���WjP���_�΋T6h��칈<�>�w-�R�0@�Gv����h{�*a��	}ۀӶ����c�@Oנ�Zma�;�y��zy8�M|�4&3)��)M���:r�=U
s�p��Z&)ǯ����=�]�W�@i��-)��D����q"�},�xC��;��p֣������p����,��9ve��M���6�m�j��8� .A�^ST�-YN ����o��]=�=��43[�s-g4,���R�3��Z��{JƋ�(R�h��zؼ��A3���\q�ĊfS���Tdj�/.'|���_P�`�9�3���4��`N!�Y�M�8�.G�E���N���IO�l��fgɻ`g,�;x?4���l�!�F�B�u*;y�o|@Dk�����]*�n���	w��=2�n�͆��,�B�aP,����( ��P|J�v�boz�ec�n�h�����-p(VJ�%�u��G�,�Q��'��--�q_f=/��c�#���q�>ӝ���}���5�?�;����r(P؅��V`�r�K�$�C�<��w,���v¶� !T���R�������հ�}���=WdC�F�]r^���#}�Ӎ
z^%�@��,K����d	Z�/�{R���|�Ph�ր����)�6�xE �@��2Y�(�l�2PV�Ŗ�����z8i��n S��LC����`��*ٻ����\� 6�%MO���^h�[��H4(�¾f��U��u�D8UB*��XG'|T�tv���U 3��Z��(i���ם�� ���b=�8��C���h�<Z(!����>_��#�m�\��LH%fX	�*;i��*����9���q�oÔ�N�N�sҢ��kE��o&��t�v��/��2�f��k���T�S�켎*����([D�Έ��T�����Z��(�l��C�������9��[�ʁ[�ټa���BîI�p�Uj�?�?c+O�K�u9�c�����ЉA\)�p��u������ǵR��Tpo͊'������ �j����G�)���i�%Fp���]�_�y�<JlO3��9Kʞ���y��_G'�++^��m�lQ�K�oMF�f�5��O��TD����ZR�F��f|$�)ω9��;XTc玥�1�(a1�gs������D1
�o�Y���ϻ���+T�䇭旚���e�P�$&D��� �׌�߽ztrz���@��L}9嘔��wI��B����7j���T�f�(��"rU���i��f��P�Ȩ�3�'[��1�W��_b���C$���G���u�:�4�|�DYa��io�8��J0zd���������Ohh��F�.˳J�l.��a&���T$O��n�u���0^�dE7���\N�Ҿ.�0t������S��rB�]��j���A���D���ݾ�6%ផ�h��½��I��iC*�};�?G���Ft2h��Q�g�yX@gk��H?A�������}�϶Ͼ����ʨXFP8ʑqvo{c�n�<J�T���J��x*n�@�Z���a'+�r�ir/"��5��|^��W㬛Vw�3�Uh{8~k/.�t9V��S��2g�d�=��)e�d@��r Z��h\��:$��T��UԼJ��b#�TRJ���Σg��ID�:��oL\<B�^����,�_W��={C�����)b�����u�4|��/�X�]�ؤ��H�M��b��{v���pp̶�j�\U�5�e8�.lX�H+�8x�Ⓦ��ś���!�R~��z]�K��o�+� |�b�{��ˎ�z> �Ǥ����#;|�1��XA��0�>���	��q��wz����ۙK�M� �u|^Zy�n�9o�ږGa�� � ({8Sg[�p�Su#���k�e�r�@ƾ�#|��PyZ��������'� �\WŸ�A����!�j*w3#�ǿՁ�0�1��el�_ewF�b+:�(�5,�.��hC�H8�u���/���Pu<�9�6��5x�߅��!n�~S7G�C;qۣ�����'���Bs���I�U]?uX�,MG��Z�=Z��@ڃ:i7�`�s|�NQ���P��Q,o��>���+]M�q��պ�=ݿ�y�#��,K�-t�$��"�)6��?I^�ʕ�Y.E�eV���s}��P�B��+�He�� ��:
�T!ϊ���=V�Z#�ʝ}�rd�3K��|߶����W�v��#��ڊ8yU�){�:,c�w^4��a����N�2˗�;æG=��.@���i��Nz����{ޢ�6�f�4L��Җ��V��_��Ù~,*��dv����o�z@�)T\�!�A,p\L�I/������~Ɲ��Q�OG��떦J�h���B��iZi
��Hl�!d+$�Y�~2rGԌ���8��lK����Pꘋt/�KQ���J����hq�8κ~��(iU�p�	�.[k�G5|�~�WϽ�X����ҙ�B���.:ɴJ��v ���c%Xj��}c$X��ꨟkJa!�Lv��P=ƞ�p��~��r�+A��[@�,TM�c.)�o��cu�Ea.F#`�qU��e��v��_�4�:8�ǣje���T���ػ�ӹ�A����YmT؝���@\2�e���tg%ix��<�kyM�Ƕ����I�(E=�f�' N��#�}�n|��6�lQl��`�16<r�kB����W�O�8��|{���(��o����SG"���w�{bo�K9|`�pvxj�g�8V�����4	l�X�U������}�+���l>��ҥ�DR52o��Z�{"����d�M��;��x+��G������٣�{F���i"J��T���d'�>o��9��DkS�RD��~�I���jdrdꨢ4�O�&[俀��� ;K�tX��ND�<���G�]��t;�/����+o��qR��7�g�j���4F=vߝ��XH6	;8ҟ	{Ӏ��OB̓k��[JP���(B1�ق S[�:����c����V�����-��$Q�gź42jZv�.�-B{�Q6�+@�0mq����2WE-��h���\ �&~E |�5�q�����>З|��y�Pdo��'fĴo7�]���bb��M�lÇ�X7��V?��T�$�n��-���jr�0�!?��{�?+y������ݤ�� 5�U�>�U�c3�x$�4~~hk��yJ�W�a�&��q����>vA�����_�P^,o�j�<�Y�#桍`!4�?V��� ���A]�v�����|�j�w0Ӹ�Eoԃ�����Ô���h
���'�\Sb����:��\���+"� nӱ�v��._��\�J櫩���q� ��,Մ�4!��������l�l�����e� ^����'���9������
e�"C�����<)�!k0t��1�<���ϖ���nKT����1b��>1���i�A��r_
�btvg�~(�~Ĕ�a�+WP:��^�ķ���;C2��aƤ��_	\+�-�Zm#˫�d�Ѓ���ύ|����5L�X&��#��O�^XâKB^7ܘDԉ���z8�Ĩ�z�>�B�;��D3���g�.G�u��*	����О���x��V�-�;$s�2	�$�(N#�t�o'
�����V�����uD�P�����}��d�!���e�bƄ�Y�6��N����'����Ψ.���왤*|�v�����/�1��H]�hbv�8���b����#L�_�|�^cM&(��bŢ��de���cV�	���J������^�Z\��w�vIɘ�.ki�T!?�#;ߓ[�{(��T���Go��EmAxf	���'24~����q�ua�ȟ��ihl����h�"`Xl@nvx��F�D��1���漅�E��"��P�~�M���3(�j{��L�*5gS�G�ä�A?�f�5�����'��x�cs��#d��g��s�AC��W�/�#o��{Zo	��U����]��mN�	o:���T��l�d.����"�����K�D?3�e���a2Eږ�/�#��u�]	/yh��E�ok�Ǻy��<�*�͂Su�s�T��q��\�w���m�k�@�y���H�[NNS��^V����ΐy ��؟{�uO�9X)���ki�2E�]|ӝ4%�&��~���	ӓ��X ����q�0�y`z���s�0d���+���)�oO�/�� ���v��W��5�3Pi���o6v�̪���
�ލ4�*����	4��]�Tdr�A``�XD���m�;�(In @�rⷑ����m<�� rټ�8CH�ü�[$���e ���q�����8�B��]/�#�-�A�5���>�K�����!*h��?gΔ@�uI����"��`�``R+�f��X^����Po��Ȥ�cư\S�ȾXW��L�z�Va��ԣ>���~��.����Կ@y�	�k����X�_ |�}�?r=O#'�)����$#�+��=B��4R���g�͓E��p|((dn���t�#��%݋#By�wh����ՃT��+��m�omq�E�2bC���W�:�0�o�\Ѹf9۰!�z��5�@���WNb�-e|\���KodW���!�ğqOq���ᚰt�q�yEo�2VP���}�������%�i-���3f���S$�%m�=�䙉���za6�,�JJ�|bm�^��bԴ���[� vYv�c�?[A�\L!��ǒ�mk=B�Sjƽ��OP�$�$~�D]W�d�)*�_�hȲ)������˚��������LGB0oH&d�콪����7	���>'�u����$�<��Ò�v�a�CL�%�/`߮C���1�2�
��|&^��>�Rn���*�[�!gM������i*��)[�1��+⌻!Du�:��$�V�u�Z�C��0��1��5���q#��0�F7E���%g4/�^���ź�	W��ad��y�P�BZ������鬥�H��&nr` ��
�M&�%G���wh7� �	��?�o�**����p��zX�-�� 	1UKjs a��j�Nr)��ek�s/��.�b�7���c����꿖�ts��Z|�F�\ U�\p���&�:۬��&�b�z�5�Z�X�_��z!C��!#��SlZ���Vg�=��Ay��Vi�j��Ze�V�O�ɹ���ya��g�Ye��TV(��oe�V�������QZ��������i|2|:7���M����P����ID4��'pK���e���c��)����>p��`����C��El(�P��,P�����W���L-��zYOG��N���!�������\v�Un�Y��~t�S���N����Y�C<�̈́ ���QJ7)���I_����3z7N!��h&���&�Ӥ���0�5�L�� � ���t���������=Y�-,��� 9�������r!ԇ�½N� �
��1������$�TIH�n�7��d&�`r,�/N`�D<X"Mb�f����l���1ŝq�Ft����VWĆ�z.Rb�Ԍ&�{�wڣ�tQ����r��^q��녴B�j���'���C������S�þ���P�ġX��`�m�X���$8aܱr!�J�Kz!4}����_K�� �����[I6P���;!G6�u�i�x&��
��"�<Oߡ�F��g��y�0�8]Q=��M0Y��@D{��2 r7�DnԮ��J���z�k|Z��sχ �l+�ɷEN�0���E��:U�{ƪ�³Ƞ����OC4]�O~Va:�U0K��8�na���R�?	́��Rw���eY<�|�<)Ӗ����l�����BĠ�cE1��Љ#���H�ң�V�tϳ��|�7F�V~�i�l�>�q��'w���ZZ���Ű �6<I�^�J����59ZG� � ����!�a��EAMv_�$�"�ػl�����WC֬Qr�b�G����GK$!W��ǃC�������Ȱ��rdr7���Dt�ӅK����������w`�#����\Y��X����
�q��O���{av��`4<b]nJ���X��dJ% �Yb�5Em��<�e{(G@p�e"�M��Ac��� &�_��j.q��8n�
\�8��d]���H��K���e�2���b�B0�θ���J�/�n���:L���	k�)����9N�Ӂ���%�1%Qv�����jq��8t��)��ӕb[	�'ސ�Ƽ$˛�b�\��u���d�5Ǻu��gr��O'���b��f�(�����+1�-L����Kr�lɱp� �W�Ƌs.!�m��
�G�]�Ǵƀ�-�ZO�r���ʡ!����3��oXk,,�?/��*4�.�t�M򎃞��HX!���Sfl��u�Wz�������� <��ﻟ젉����� �J�T�(��
6���^�<��M�{*V�uԴ|����]l�e���׊^<��!,��w�^� ��G_���숿ͩIS�dC>��2��|is���)�d�{?mm?�dd�m�?]]��X�zKa`KSJ���<rAa�r����?��Q ��"�`��+YR[.��aG��<)?��bX2���#���!�G�6"$
~��A�-r�����
��=��E���;�� :�R������Đy��ox#)�n��Կ蚺#w�XOF%zmU�9��/���s��:��b��g�Y��ee�G��?��d2�;Ь�������V��K����e��(]�U�:4;�%sl|D��u��[���u�����%GL˜��!�Ip���8��p�]���������R��1Ȯ�e�B�ז�CQ���;q����z�^�"��,�c5(����1n�u��){x��)�a��7�8�F�a��mY[���� ��yΐVR%��0�k�XF�r�_\N��!�v_Q�)�*�S1�,%9M����r�W����Uh�&^uHA��fqR�if��8��	����b��NW���M��@y���F�qsI�ҡ�%fJ+�Y�Ma�A� 2��6mO�k�j����,5�D��+�݊�}.���a��=�aepImf���t�%tsT�hwH���r��_V)�[&8>R@E~?�ʲi�� ~�� �d�y-��:�����o�H=1��	��?]��������&�=� TË��@�a-����"���D�D,���-�C�_A��R��� !K�R7;�!ПU�u�m*�W�*`�O�5�:?ߩ���3�JDԫEX�ݕ^�ki�H� �|��ǋ�)C%jSn�D��\���-�m�ij�&��ʈ��a{aĳ�Tn�?���"���(^��O�j�@��G�� wRc������ȭ{�R������c��a�4-���!h-�X�f�iù�i�
trk��*�FqY~�2�_m>�"�6M�~���>q��6�k$�\SQdD��_��(�C���b�Xh;D��'0�*���X�P��0_RQz.##r1l֧�x|��2'{��*�\��<�:0����D�B2�"�"��sߘx�hS�5�kE�̾J��Q��*)�361>��e'��r3f���op���a���{�ڮkr��^��ux�k�9�m��.�޷�p����:/�׌Q>�����-A0&������n䆒ˊ��8P	���\Ua���F�	8���}���N!t�,��R4�}:��
d-0��gk�Q�i�g=I��݈�L�9�t�CA�d�6ϩ�}"r���҅�ĸm/�AC@ro&�1����_CZN�ڋ�+%.�L�)��E��x\"G��9�L%�qY/T�a�ѷ�͛'��3[Q����K� ��|�hq��4E�u̶��M».F�j*�uP� �ϓ׆���.��`�FJ*}�d��K�]nE����p�����i$��Q����R����1MD��?�,>蒦1�{0�������5m/��p��{��Y��ɸ�2������7S�����$�#L��el�rc]{��=�Vz�'����}�b	�B��P�\�̈́_* �,�R�{�$ٵ�,��<�6�ԏ:�6Z���`��� ?�j�$��[a�ou��S���WH͏d>��X����+na�ˇ���:�l"\��8|�Ր���Ƀ�H/�6Z�Y�[#���'�!d���m�љy��҇㈢Y�}q�=\4b�Aw/:.#d%�L�J*���U�.ol1_���7�E��(v�>��,��v-nR�f6#��UwG�V酋�`W��C�<��}�vmb���Q�ƨ�S���?�@���m�����Q����<���Rߌ(C�;U�bJ)�NJ�m&3'{Z3�g&w]�R�KD�K�ݜ��Y��tϢŬo@��I�T��i�m �S|@z��x�7��F�a��A��̵<����+_S����B���� ����;���&�'Ȗf�+���~� �q5�8���� �f���ف>0[��@��K�T�b`Z�@��و�`�v�ubnL�Rw�g*}ʫ|
��f��5#��P^!J#���t�j�+����	��N���͘�<"�W��
�#W�%'�@��j�Xfd��|\ϧx]z���??�b�5qr+J��`q�ԎD�ä�J�e��y��?��^�����C�+P�	ۻ��,�Z~��Z�s)�x���]'HUD��%p�>���}w%Mk�lZ��?a��a��e�@��J%�z%���DGk��R\���8U%ϧ'x�� �i,�b���H���|�_�ۣF:��u�5"4���+&����e����5��~>��,)	;2�/T!ˎ�>�
$��$a��gF"`i��'Xw�E4.�	o2��R±�$��p��.�AR �7�?+�3������hC갣���<���\�F�w�n����V��B�tQv��g٠sD��o���ð\�Y�	?$œ�����5�u|��Q	�2��vL%�u���Lת��xl�z�"O7�]�9�����j$��kw��"YUU��v�9No.9p�43���1k�̦*Ʋ���SR�m���θ�����$U3!E��{V�w�b
�5�L7,�޺�K}�2��`!��3���>CC\�E��D���2@�~�$�����0�;tP�8�
��@C,�n�ʮ^q�7$(b����4�$鳍KL�ge���̹ϱt�����V����F�/Q@�w����eS��ptD~*&��#� e�nյ��>�,�&�f����	����ʫnn��&1ٝ���mPh��^(=K�/B '�`ĉp�ʪ��Q��x�P �[)�B�t�@<,{�ÄΊ��P-�I��tM��w��OZ�D�[�W;;Y�1\&�W���*r_R�'��}5u_\;�#Wl��mkRM
[Q����"J ѷ�Q��ė�+�ܤ��?]v��m�|Ԑ�5�P�z��ʟU�HPM9����5] N�ׂu#�(�A4���ղ�oBv�-M���V<��Z�<��b����Ǿ���JFL瑶�γϦ�
�wWp����C��!ם��`⍐f��H��2 ��}X1����)��4�M�z=WB�2w�~��"��lV	t�bS��&0��\R�*e�uZ�Bt�.���˟uK��6꣖��]/Zc֏<���G@Ļ�>mAgM�����P��~��5(��gi�0j�x2{%KN`,�6r���d~�gR�F���ރl��Cu�" ��֐�P��aU7���ˑ��EG�q����OXU�$�q��N�&��5�c�};�mT|�e����9�����+���8d�����o�H[2N`�	j�� �;�J��ɒwG�#�Q��f��X{ԫ4��q��V{�-
�]iN?50x}�i/s	7}��@���P�8���Щ^�|$L
��E��fh���/����*�a�F���y��n�XDM�?O���ˣ�f����m����Sxy�	�D0<�/D<4�s>�'�A�֡��zH�I�d�ۀ�t/��;4�9B0���Jr]pr��vp���$#�;�~}��-�є�c�"�2�֩ԉ�v)�bɡ�T��,?��ĸ.�M���IP#�I`�l�R�hξ�A��L�{G�I��p���՚�h�j�?�>(�n������/�H���keq�4�j��?ˑ��c!�(X����{'�,i�WC�oF3�k���=���=z�U�K���m��}�1���$OMg�B�PCC�Q֢Ԅ������1��'��%	���:$����r*�8�i��5����p���*p��'���l[���u$���T���N�D���p�^[ T��`{+:��m��r�P�y�>�$�݂ƈ� Q�����kſ6ɣbckU�����ch2�}���s�:�_K��-%d���Knq*,�y%6%���M3��inx�mΡ{��>��>��M�Lf"&�#�i�JXI+9n�B�CB���q��3�oQ�l��9]}*�gQ
��d^�&S��ɓ���:�
X&.�MK��y5�E�N�9�l�OL�Exbi`�%ۃt@h.$�o{���+��J��-��������U:�u�����C����o�ը7�~�En��u�f�q��;��Σ�׭��#���n�ր+��O�c��*c��6@�s]S�[��_�Y8�A��${��u@�eG�Ԍ�~Mr�ѳu$@��yT��L��Ю��j �_��D&��[1��<���4�E⩊�y@�&_b��4'��N6ʏ*����;~��#�P�=��7G���Y���:�T�����b'�[KL�7�狤���0Νd��z�>�$t,w<�[ �/;GWR�$i�d]<%p�y�|�����Q��DKz�"����K������,��oc����`AU_:At���#�H�`�t������Z'�d��M+��}G�zg���j�~�	�����i-S���Z2��w���?�v��א1]��lS�����Cw�X����rk��n���Q�}��JM��v��i��kLjR�WT���ù��|5���'���lu�w{v�bk���.��
�O��Ģ}��q+���1�c�=1��~���1������l��]<c�����5�>P>���m���D�;�q4�O��X�WE�i����x�=Pp��:��'���mJ�z���6Fq�5�$�02��w�>��<��),]U��Xr�.g�C#wJ�8�(����C�xl+�]_�}?��)R����^�d��(�-����B�!y�7I�X�TC�0��-]�P|u@����"{�'���)!TS؏{P��f�5�j{��}o%]�,B-!�뗥��q*v&l(E�B���7�7[�6T	N�]�A{�������Z��(� (�+圩�����A����nk�B��LFr����o�E2�ZTW�VZ����+l�����t��&�ah�U�L�s��m��=��e��Y�tՓhQ~A��#,�5�J�	u�+뽉[�v:[��̂I��1i�<n�m�����uʈ~j��6.h]��Fv��u�����{�"�GjQ1�Z��J�����:q%��q�����G5&}�cS���u�0��wŸu��䡔�T�8�]qA��-����ö����0G��9�L�D�����Qڨ�;�zhR�����ܩX[�p $H�05�Lo�9/�]	 Q<��R>�&y�'�?#�]#X��}�k*�o��D�Ȉѷ-#�ZIj�vEdi�ˑѭ��M�x������WX�ʢ�������qC=����óo�qI\;=�*�i^aW:
��IYa���D�(�	oRả�4o�M�w�q���W�����$Æ'�X"D��EP ��O�܄j�C���G�̈́^Tu��c0��&���Kp����
!lK Y`��L)3��a�L�JΝ���=�I�x`ь�d�c���6�OrP��c������U�{�լ"�@t��!��C~��3�NЩ7���y�e�in�J3@���hїߓn�"���s]/2p`�Q�)*1����)A�����OH	�d�gc^�l�L��-��`|��v:��ID��-���q\ؒ2�QLt��������Z�!G>��
���t�V���xBL�ʕ�/'���-䝸F���1��*��{!��v1k�UD��CE�`ݤ$�0{����ـ p͝���,��&�/2U^y���˚�:/��h����z"��j,ZW���<dľH��=(>�:W���(ТJp�1-MbYv&Xa1�w(n��}S5Ĭ̘�\��
��b#0р����62*���O�Ou(�Ԁz�Q��o�N���i���� ��"�b�����J2=�X�c���	] &I �-��ޝj5�ܸ_�Db3�*�\�˅+(�m��[1B���;�1y�"K[���pw���R$v��p秚���p�bW��k;uժ���ﹳ�����m�����VGb��'1��<�rX�B�� �>���#�:�ĿI]�J#�;�l{b�jI3���k�S�o���`ys+6�l�xA�P�0��+��u�9� ����a�ћ(p��|����wS��vx��V��$N��zO��peΑ��B#�M�D��'��ŭ��;~�(سr8�T��d�_$��V��#Se��*,�-!��$��
��{��0C��x�2�2��c$i���W����K"��#�������a���A���o��L� P�G)�g�|�q���>�O(hQ��Te<f�LN��삤�?�>	���J�}�x�ZX��(���zf�t�A[��ko���r$>�� ;��P��4L���vk�W�}g͛���8h=�á��/Q���h�E=\�� :Z#�3�-}��V�	/�S2h��;
��%~p��}p���f�{O����M gf��m��	(cY��4���lj���9~B��ź�1E��.~#g3ث#mF>3�K3�=X2�D����Kg��F�^c�~/��4 �g� �T�ʃ���
�R�o�w��,��W�h�ĕ��&�Zn
�9Js���x3�{6��\C�S�>�u���\T%�/�����0���A{��X�+n���3F�/���0A�j������]j-��p��A>�Ұ�~�@���@�O$Y�����n�4t����L�7΁�v��5�պΛ��<D�>�{JCo�|u|�n/|�&K�����$Ǳ�K}�|{.<6J�[�������I9JP�9y���
�=���JǏU^����������$H���!Ay_��6��4\���8цt�||N�t��G�ƚ��k�I�������hD�28�2�I,J	DY�Hԁ��(�'��W��\��dH�� �͸V�f���	O���P?�8�:d!xƋ��d�B��'#�c��!R-�j�Ny�	�,�J��/Vk�-�	��)3��=Ȓ��-������|����]I�7Ng���`��/��T�G9��X$�6}&W�����MG�I��>��Ö(��)��z�~�O��w2d�]��������p�k}�_dY��e�_��=]Zw��6Y�� "}���7�B4r�{bm�0���A��	V�7>�y��՘�F������ [^(��W��u���(����Q�������N�	�N� <|��R�S8�������O�p�
[ ��}�<'�82��zG�Q7��}�?��L�������)V���T���l�����=��x19�����>�o4�dy� 3��͞9.z�ME�.��x�b����F��v�oTB�������(*:���K[��3�OV�&���L�}��W<n�!2d�A�_{�����9Bf8;T2�:'��x4��`a�[-~g��*�\>m��- Ѧ�<Ј���Uouj�Qy�`�ד
a	�r
i��]�r(���?xg�L^VϤD�ɥ�4LD���d�S�.)<������D�d-��[���)q|��Њ��C0t��l`�ӕ�u�ᰐS� oTk���R%�R�X�[I`���.�8Q�LU�j��#���Ƅb#�d��H�3<v�~i�,g�)�<�W��PE�jq��Yap�p(���w�X���c�D9%�*�ox	���O�6���_5	ђ��C���������С�������L���n]��#
�/F�O4�s�B�6ۚ�G��Br�}��P:I��JH�0��U6k/��Mh|����D }O��%	�CM������Wc1���$>��N�ni?m�.CB3+���ͭ��4��mP�[:��}~�9��W��+s'h#�䎉WI/�v�`��l�'��MŐي��_���9�s��mI<���2�;|�! ��[�r�}(�u^B�Dw���푂���M5���;�JAr�+k�g�{KMD_����Se�6�)�T���N�|Ăv��0j����2,z���8U�	B�G�J��=b1�'���׳�G��.Р?A���-澭8����9�J-�]��ľ��6Rg�}��A��1Zp��%�G���*aN����'���g8d޸�|3H�uc(l݃*���kYv���THK�����M���ٷ�D�v˲2��OB���X��k��nLE�,̠��&h��l�X�����0�p9���Q�˒٪d�"12��`�B�)Á����Eam�iA�{;�:��D��\�.n�4��v�һ���[���\���(w����s�8,�U(�DB�_i֛(���a�n�Ꙇ��(��(�-T�؀(���ɢ]��\�C��?���s�] �*�썔1�.�i�B�6V��t���U�^��$��y��m-���pO�9q@Ӕ��S��z~VD�a^���fp���lO&�K�y�� N���v���o������h|�P}IB;)@�6�w��#;5.�
BJ�,�΍!����_�T ̭Ó��}��ۓ���%K?��mj�t��ͧ�s�:�ݑk{�Z=��wpG�˗1���մ>�n_E�_�g�6�>joq��&��L`<}a�DM9,���g��Uv�7�Svm�.��줹'(.��put��JV����J&�ss!�������eU[�
u?��W9 ��$�,�.
���ʡ}�1�<��8T�5�3�%�,S�ёŻ����o�=��J���2O9_����+��Mk 9��w��Oat?��G����{M��f)'�p������0��A��|9W��n�{0��=�'�ytFϭ�8p�� u�f�G�1�T� �ٞkYF������`^_��&��k������I��q���=��7T�n�a˳�B֋���{T�>"��s5=L
w���e���D�Y��Z��oz�6��L�����:�u�1Lf��͊~���M��̇���]��;��g���]��4����2�$�~rIp�-#�ŹK>�\'�n�B��d��K8Usu4��B�*
2G� ��8vپ��pX/G�~��].�����|�a���P�6?���d�_�����A��C��>�o�
&t���@����E�Yn8N[�P��?�w<��f��d�L9MU6[0�ZE�@�ͨ��k��G�Q�
*��-��Y�Ȧ��L�O���p�j���0�Ǆ�ݽ㓺Js�����8y؎���V���}q��UU$���.�\���at���-�؄)k�'܃�^��d�4��b23�
��R݇T6!�0�eh�K�������G�����Y�kF��FIpΥ˧Xr�3#X=q������<�^dm���f1��T��J	�2.Ck���Ë��O�4����
z���ݹ���ہ(�?��
]�t@�%�Թf�k��aϪ�M��0L\�!����D������r���_��w�������y�{ �T+�J��U�M�*u@|� ̾v��}l�ǚ5o�I��q�7.��t�sn�ve��Ȫܤ~�{��t�^��)�G��Uy�f�O5wu|���g!�!��0Z�
���KP�SO�'�>�
t~�s�(��x�.?�c�&`�p�!�^��~���K 7R��Z
��-�\m�|^ƇA�l���O.]L�I%Z�<y�5^P���qG�ן�!v�;n��2Q���ۭ��/�
NYݠ� 8|R��I�qA{�t��Š���U�.4�~����L|�����)�T(8��N���gfA�+��#��k��׀}�T_f��b��P` ����~U��Q���M�hذ�����v�oO��P�}�V�7$Aᾞz7 �/��(	���s����)^PC��b��.7)hM/�YJ����m�> ���tU|C�>y�x9GT��o���χ_Ѱ��C�D�a2��S������X��X����~X
Bh6���d�MV��'o6���x�#韥�	a�e4��]�J�k��&���+
�y��9�j��y��(bjG�\�6�(�̩v}0�^;����hcdK{��B3��$�.��Q���܀���.h��&$B����Kh��s�3ٌW�2Y7������~�c��fЩ@��~9�rZ���H=�E0	ؑ3���9��0l����F&Y?!]8i���B�JC+yZ�gɼc�c���V�O)��	胢/eξ���[��x�O�J�6
Ռ����C%�#�[����=N��O�$��G��iN_�	\��|���O	�?F�%��\��Ǖ��Q��\�v˯u���������(�F{��8���Gأ	Ŝg)��gg#�&�����w������=�����`m�����pE��/Rzbܙ����V:!��Ȳ�d*b�v
u����(&p���p��/�5��%�o�	�X2ê)�����_��S����\��)ߥ�ϡl��W?���5����F����(_�_�1�����7���A&���>�^j������n�Y&G��ɐy��)��
��T��	W��iO��o)`�n_n��GE�=H�r�]�3��f��3��6�(�-���!�v&��~��W)B���h�!r}�LEuSA^�9���K?: ������F�Q��0`��5[��N7���v��ʥ ���tv�0�?Xߜ���z�(r5;���>��r�����D��_J�yɹ����/{�|������B��o�ø7���ό�Y��5]��<��t$��q�n���"���8�[��3��#�lab�%�����?9�ȫ9�&M��IV��������[���*��OL�/r�}�:�0_��nZS��r��zW�A�i8Wq:,�'�ଘ��~��0�B	i� s/���`�~֠����K�<z�K�!�ԼJ�Ǭ=��[�iQ�Z?�S(�ߟڭ,M�޽��^7��<8Z{2i�b�OMM���c�2ݬر��5��;��"%D
��^K�H���U��C�������N�Pk����
$���C�
�����V2Y�!�|Z�k�AR�<W�:�Ơ�\GE�AR�3������eݫ���@�W�o�^m�;����<+l2�9��2?��
�蹕lL�M������4���E@�cN����WCD9:�H6�0o��7�:�?`��|�`	5In%[x�d���Q�ؚS���bp��mr�"�n 2����_�k�<+�c���[ҹ��R�\
���Fe{���*U�ݏ�}�ǧ����M�V�wxM���a~\����*���T��	�y~p�;)���x?A����÷��u�ƾ�/�i2w���g��i3�wS��gE����x��$"��Z7���8�[�ϟX{M�wN�JA*��#�\^����C �wewE�I�Y�5�/8 T�UGYs^�mk`N�����Oˌ�z.�e{�����G�ú;��r����
��4'�{Vn��Jq�9%Z���||�^��ķ�7
�8��-(�GF�3<�'<�]���z>O���L�$��D����[SM�ܴZ1� '���l_j@��s^��t���+d&�	U�$a1O��#C��S1���F�T�G��W韺N���9L<�sRp���&�Ʈ.��3�}��޲Y{|����8�\��ײ� ����|��+'��qXDT-W�D(��gN�Y%�b�U�"X&H�3���e4q�d`Dʵ���l̩��J:�[x����Φ�S�jQV�K"�s�� �?e�^4��JZŰM&Ҝ ��=+��$������4+��iB|dy6#S|5uˢA��s������	���;_�#>�&�0���v�����6מ� a��$��22��U?m	��g�~�mZCnCc���QQ���%��j��͔MZ��K�5I�.M�}�0�8�m��LyE����3c�Qn��3��1�I>埄�7{��$��R{��g�d�Y��,�v�����hFD�_�M0�W�H�Rnjc�
��i�$�w���!�	f�U��mьL~y��W ���ι;����������L:�X�{G`DD�b�B%5���JO9 B�=�ey���'���&����%"��V�UG�Y�:���F;���	c��	x��OC��k�Q��\Zg�C�gOb'N�+��oBܙ��������j/�����H���E�����f j��^���Wii���/�}�n�Wh�Frmf��V`�sսBu�����&�惽[��X�s��u��uԮ���a��{�ƹ��p?���*|(��Њ#mi����3�۱��.�	�[�E�h�$�%�f�q��V�	Ŵ�p���,o(���%Z��}^��z��S3�&���s9�[������LV�QKͫ���"C��gb0f�#��!�u�借o�k�0�*NX7�U5��3^�XF�j��������$�Ւ�q��/P���o�ze�K�߫��?�X�mw�_�T���q}�y.�6�λ��htH���K@��d1�cXY�s@�?l��^T�7��]�
���W�/��LG��^�+��|��i��m��As�	}��\��u�!w/'-��i�VN��Ò�sI����^����Ђ�gH�&�?j�J1�1l4.�S7���۠i %�0�t�H����IѶ_�$�Sғ͆���60싨�]��2[%�e�W̚��rd��н~����T��pV�3��x����D�Q���="�����+5)?�7>���{���3��z�z)hbN!�" �s���/�k�j/�y�%�����M%2ж��c֯x�5���ec�s�=����f��/7���;���`�I$�[�ҟ���@vz��h�r�A�M���;�=Q�qG��/�p!�Bb5<�ۚ���1�˚k�ʚ���Y���|p6��^�Ȍ``I���oyUƉm#k�G]�4����O����K�|�~	Y�)H�-i�ٿvX��q�d|f�]�f��£��ӣ��>�s��#��u�,�dB�"3׽Z@;�rh�[�@��lZ���:����p%Կ��c���f�VO��`KP4�BX���~��wI=K�y�|e��+"�a��� z:�`��c�L��RԖ�
�z�He�G�s�/H���W�N��i�4ܞ3�ʽ�a�3r�n.�j����l�/"�v���K�wk��YDoȢ|�Ә�C*�}Q_# ���@�v�Ay�a�V�-�.6�g�/<k����'7��xMK�k��
�	���h���<�fk��k�N�;����qF�&t�ai�]Zۮy�
�_����3Nj|ae�̞��m�[N�u��%�9%>:�+D&��R���G'��r�3 h����I��\|\�o�z!*ZYN��q�^&���H�8��k�6�q#{ِ;C��T��΍T6jw�!�9�D\GN��?[��g�
��Un�{�Y2�k�P:�ښ���d�9�!�B}l�&��
���݃��1��Nl]�ʶy����`S����4��n�q��Ёy��4y0���#J�1X�������Q .��(Q��Ӗ����)^i_/��oT�}��\�����u�H�yp�Q��*�w�`��o�X�6�j��t�>�������&��l�5��n1.��N.�؆^����SoȚ[��U�;0�o��d���%[����e�|�$p?�G�q���2ݍ�nė�S5�4D��@�F�%�'J���w��#e��$[í�QO��ƅZa����@�3d��Xad�'CawAZ(�zJ `����B
��f���� Cup��	~�N�@ݯ�v�><��~��R:.�߁QK���\�L���P֑:T�IM` ������`fT|pHzx������ ݡR}�ᘨ���cX���U�V��b˫�6J�v
��5��P��P;�B
�_:�Dt�����4����D�2�U�J;�ͼz��K?7e��zK^b>G�ߍ?�q�ǘ��_베�o���1�����G
��>e�#��!�2g�\���u��+Q�����<���!�ȿ�ݞ�s���l�U`_D֬�% �`P�m�,rp��8�-O�W�9!��f�4�p-V��7N�ĉ��M Gj:��_�
=	
��4�F��G?���	���ޥV�I��u���Tc������QP�J�Tv���q��9"�m��8a�U������E�̜E"�0cv����l/*�������aڦ���nQ��;M����2}�5c�K�_
-���@�w�̳�b�)J\�RA�|�(m�����QyX}�0Q/؛抵+b��ׄ���V�I���gv�^ru4���3J�/��Ҹ���).!!m����'��*L�s3x���d�O�恽�!�V��;�XZ\ ���'���P.����(��.'���"m+��'�/P8P�e��D�sX#����7cY�p��X��ْ�0թ�F2&)Ch���r(cHv*ϙ�T;�e�JM�~^�Do��������4�K��\��f����	��"b���j�{:ZpuE��8��J���`xۦ
E��I��*EB�J.t�>���A�M<~���ڜ�=82�F1��!�P��Rī�l5%h��g��	t/Ӊ5��0_�&D9|E0�&S%4�Z��l��`妕�in�� ������N��gzrP=
��\��M�R)��>���h��A���ďA6q�n�����.���Z�',L;��4m���NT9�(s(��e��%�c�H�򚡫�Q����JP���G�.�汩ob ,��n��U���K��<@x]������F�����i��>I�w�"��F� PO�x0za;�G����~Gc̣�o@�,1��~5����������UU��v�� K�#��!���F��˦������j�'o�>�!p`���XGu ��l;�V�4�M�|ֺ�ѱz�X�����Y:��.��ڠ���ʵ��ϹQ1�Y��g��aY�rdt0�L3L�@u�+�Y�����[;���H�Aܑq"���� ��iY����x��<���f��ˑ��i��>+�1%�p��B{�|2��\��M�5]S�Ўĝ�_@E�0��\�摦�&}א�T"v-�%���x;�W�}�I�ta���(��e��7O�� �%\��*���!�?�qڀ�����rC��K.��^���ax�h�#[Y��ü����Ms8Pr�|Og� ��-�8�;�m���J�ޒ�?�|��W�H��t������ضޛ�ڠ� ���v�}i�O�i�29Y'ۥ7������u��.^�����o�'@ji~��Q�Q.X���n���$���~|(]R����jW@�9
�Wjp�O�����4�'e�h��:�������ę�fd��?���_.3��y���"��bW���藇�6S��0)x.�'B�X	�n/���W�U��j��j�YK:KO�gu"��3O�$�.5�K�Ktڿ���o{�:���<���_�BC�P!
)���K�x�%Z� �Bx_�N���;�o�j�Ľs��Us���D�-��TN����YZ�{ݓ��Z+:���>PLF�<��a�#��r����E���E�<�W-	}Y�q���X��=e������;��f����z�BJZ�glW�*��p���/�TW�8�<�3��>����f8I�.��G�S���pMA���S���d/�ڞ��p}f0_��g��MU��.d^�����B"��wO]ȱ�߄��(���L��?Y��$��hO��3t�jOUf�P��+L�hMGJ��� �g��b��lh�8ҙ?�1���yxD����Ou���=}@���cd�Iz	״�ΙTB��9���чi�\��v�C@'L��X��>l���dca�Eg�UQ� �$�7�8�����C�|]�ne�[��m7*�؇�%�~��q����>��ݏ��9k�� �[�o^r+����3ź�T~XP�ߝ��D��ޮ��qY;um�ʹ�acG�^����� �������A�?g�Rh��i��&�<4�����ц��w]�W7>Ew/p�~���d�u���?���%ݹG�Ä��_����"�,f�]����"�3Ȕ�'B����0��#�2aO�&�!��0Eu0}��A��P@�A�"i0���J�, �M�ʷy��\�����k���/uk�����o}'��s��M���DC{I�K�	��D:S-�q��X¢����K*�T'v %L]��g��E�Z���z�jM��e�%�Q���t�>�'���Lo�^�<[��@�)����-qV�{��q�2v2�q̺�1*e��"MTH�"��F�`�78���M�Me�S��B�f��Ch�dr������uX��v�<�_*E�ŵY����:��ԁ��p�^�V2¡|� ܎]��2m�ɇ�+[�݉�`��`�)����aԔ�l�������lC���BrJX������a�K`w�Y����b���gFm A 2jA�-_F*�w9[��L]G�g���ҷ��.����R��p�$�hS�
NpL�/2'��l+�S	� ��hrB��!,�}��7M؃l������>h*3
8u���|�C(�{�<B�����tXr+��ʇ)���8��趑��*���'C�d~n�,�J��Hq�n�1ZZ
�D��(k��i-O��u3N�E+�^2V�����[PnU�-g��3�s�{4��"�	��y����n���ſ������.����ّǼ�X�T���G0-3a�5 ��H���J%��`Y6�����R�':���$�T�8�E�ozV�;�����3�3�m=��_u�WOXD`f�gP��d�/�+��u	�����F�@��#%�b�������9*K3#�;�Y%>o:jo�9�gQ��]�v=̃�%4�cT-�1k��Q�#�Ma���{<g�Y�
2���X^`��_!˷�_j� $���d�J���&�M�Bm�*t~#����L�7������9RPX��=�D�f�rx�{�&;�rCd�6p�2�r�(���&,�!񂸾кg@,.�M�����Av>��[�d�����`I{��.'��ݬf�m�/)ZkH�W��\�*(����RA4e��D_(q���u]�J۵"O�Y�O���a���F�Bi%tQ�+�[���[�$���-7�>W>86ϑ�0t���g���)�7��*��TX��ԃ_d��(X�`�+��e
.]_�2�uj���r�󐨼X�S�w�������3����5{K����]W$���|Һ�����>^C����I���1bц��tLw�<�W��+_J磜y�,$�jXD�T�_T�*�ѪK�j��!�PuO ��W%;E������a>|kӱB'3K�����;������A��~p��?���i~J�?���عRԀ]�Q���_l\���s�eK*VW����K�9����>y�Q�08vo/�+�TL-&~� ���$hcʽ��a&��כ���F,M�f!M���p���]�W�7	q|�?�,kZyx���VA�;.�r�5��,\Ά�P��z'��e���j�Z��ŷ��,u�'f�0��qV�>���k��b�!��W�.�L��D�!�2g�*v��i�`�8�� ��"��LiU�i/��>��"�wX��i��qU�b�hǡ�TL�ⓨ��>O�\?�߂a�D<���Fl!�uD�����YV�+o�T�b���Ӑ�xP�r"���Ģ���^�8,��zE��	9��2͚����&4Pm@ *��G@�Ip��V�c�\��s�t��;���/}ΩH��X�4�Co��T.@Ho,ZMn[R;��+�0��F�������� A��*�B=؇�+��=L��:o���.����L"��_� �9����E�� jϔ��3)umz�2B�H��5�:�vlyI�l���#��ւ6@�HZN���DS�gK`���G��YνS4a��\eC�� E$�>̍N�#6J/�g]7��f�]Q�o�o��t��_\�,[r3�"�U$�O��%��M>�|�*P!O��Θ�܏˾g����h�%=���`��&��$҄��c��̹>�����E1�yI�w��4�������Bۚ�yLQt6>9�O�B�n=h8�=�����=8�i~���kv���F��,X�/D(�#�>S~�*a���Ĩ��lo0eܬ�������@e����:s���Va��k�K��i�C��4����E�n���@��o���0�r����:���#wq)���JeA��������~)b�ܳ�����,�W{�~���$���ɓgJB�/�(�"xqs���D�ʔ�aG�T ��M�
B=��Jx��["�mr��.7��utY�`z3���%���W���ȹA��he�G2&�X���{Y���j�w{"h�u�"��˽i�1ksu���U|�m�� �	�s.�3�z����S�?`V������\�Q��~��<���ON=C(�Ɯ�`t�:`�.�,.��3Rq�t�F�=	_ d)�bu����B�'#�L�4U����I{����
V��j�[R��r�~�+q���+�z���|E{Ϛ%cj�*0��;�i�g��o<W9�u���S	����.�on��c�����Ko�+������!��fT�\���+)Nj�
����X�@�_/����1�ɝ'h�^�b�%e�]�u����v���?o��$9�T�k�t��O�i/���c�9��X��Ң��紘�"��)m�,7*�N��D�B�,�-m���Nl}wЧ��{���_?z�|^�Ԡ&[�T2˵C+̓���F�E��.��c��� ���K���H!O���A G����1Y��6�Ć��/3zEQN��S�!Y����8�� �}��g�bͮ����9��[�%�|�������Y�7�k#�I1���j|reEN�p	W� ����3�[t�_U#M� ��k��,ɸ|V�v�X�+�Al�ԤP8'�@(85~[|i �@J���7����R'o��8u�ZU>x=�_��A횢��7o�lJĚ��r��Y�U�yuv�
7;������\��d�XaC��X��V��X�CMA[�E�~��E��'��ε�\{6k�����Dc@�P�ÿ6�٣��?���M�q��_Z�Mh�𯀴���e�g*b��G5��n���������Ub�C���7�8l�Ք���*�
!Ҍu�O����65"����o���߮�8u�R>��X������v����W+@�s�{��'��'�n_]z�|N�]�X�b7*�J*q��e�:�L���0[�W���u
�N�)d�ݜX�TTO�g�7��	�/���r��b�A�C�f��L�&ۼ���pxb�|���� ���0��Eґ(���ξ�~� ���;X��;�"��gK��{�,H㊪���t�R�y��u��ŀ��<�� ��ˣb�;�2�Q0���͈!�9�qw�3�T$�� hj>�Rݴ��y�� �&9�	�|_�<�Z���@HA�Z��ǀ;[.ז8�WX�~+p�r&�"P� ɬ� 'Ѐ8��ms��|=+R�;w4h���� V�h�Lmc8>H*�JM|�<�w,5��u��r��/RM��J�,��������ssQ�%�0G	��}{���������$�N�� ۷�3[N��+�,xT���TFq�C�n���)�Sң���v��т{�h�u�+45G��Ƭ�3�Ck,孃/�,��#$	�ҥ�k�%���D�F�n����I�?2n���m�>�C�і���*/	��o������R��8(����=n�IBg̟]=�noM��2�Ų�Ԙ�>'��W�{欦��;��f���"*�w�Yq� �%���;3�4�*�f��:C-�-�]�Y)�� �Y� Ȥ"��cK��E����]���Sbh�y��Â����?�Lt;����u���lڴpU|	ܦ����X�~4U+��7�	%A���Չ0J����X I��Kٔ��e>P>�t�wڦH5���{�4)]��Љ̅� ���3��lr��5�e��Z��EGmOm9�P�p���!���E���'�y���TM#.M��!�
���u�f�6���ħً]������w�^bE���)�>�C�QM�_-��P���I����d�1��o<ʾ��Jh���ƕ��|h��I�~���s����;�s>8V)��\>���w���/�]�7�T�P��(�k�Id����kݥ�1�����÷4M�� `���۠|uӅA��#��%J���QE¨	'���t�3�Ì��oK0��N`p,a4)�1ʳ*L����H6��B��ۜl������*�bhj#����R���)��p�a����>d ��m��Yb�W��[4�Ell�����<��q^f�%(��9;k�C�z���C�7��І��+-;�<U�rS`�NV�5	tˬ-�d�~��.�& ���+7�ᨏ�,�j?�܌��H��5Jr���������77�m�*�q�������e@�}(B
����|=����� >��h�%�!�<��N�#�y`8j�,��Y0��������G�Y��t]`�tO�۞s̥�1�u3�%ASB�H���뚣^�L3L�M|�Ls6����Ep�|�o&KU�� @Ը �)Қ�!�9�2�8�A�&��o�������6���k���Z\�
~��*L����;'�5�G�%|�)��t�@�$�2[�N�<u]�t^�q��)=����2�{����zBI'����4��?1�	��(x�M�[�'�|�:PQ�\���N5�^�Pyz<��H�RĚ�]���^wy�˯��k�w�Τ�6�&������2�t�a�A*-CZ2��Ӗ�L��nmn1�nD&\7��iV�*��[=Iys�3�+����~�A�������*Y��f�G#v�K�ɳ�n�	[d=����s�>,��:T���I p$\#ѣW���}�E��m���uD��i�E��Y�ҟ�*t@��q6����H��@�3΋��8W�y7=����<��A�JoL�,I��������,�-J DO������a�MA�#�螂?�'=Z@A���Q">wF3�5J���]5"�y������Rj\C��pj��3�ٸ׊�ɾwW����,����1[�<�?�����؋��O rd{�Ϛ��N�Ѿd�T�/������h���!��K�j #�Х
.��Z��u�}���X��v� �z'�u��F���3�4dY�*�J��[�Zኞ��DH\����9#���L�4�I���g�M�2b�pV|�N	��VNY�Œn!��_���G��O���
 �x;�QOb�2
��+�8o�2�X�>B��k�{SF�S� �\�!Q���{�
!���k��%5n7�\y܇�
b�/�XK�Ň�)D�RS�W��s�N�?������ h�����E,gS�C�f?h��{j6Vp�:Szcr�=� �5sx����߾��z!�����f_D���̏�.����w�V�􃗬�����jg��c'?�U�b����?O���Yt��^�{X�_u�J�H�����`t_Mn���\ƾ�#d�>P���2�1�]z��yR�3�J1Vˎm�=ҍr���g7�_/��,�r�F�xg�S�q�+�]��nc�scؓ.:Il��0:��`��$]�hSu���R�kyd��#�}�A������6D=��XR����)Y޵*31��@�2���V������@_b�U3?����R3����*�k+q����g����=�\�5��0�	t��{�䘯�^r�=��@e�Sd�@�5	o�_�y�^ 䖞R�o��LھQ� ��N��|�:,�"�Pn���FC�#-U�^�������R�O�����k��P�Ay9��[l���� Tb�z0ȳ�L��Jܾ��V����֬5>�÷�P8x������P�ch{�*Y~PQ��V5��}�u��,%#!8��.%�__-�����W�C%�{�A�b,kM���t��Ķ(*�!V���P�@4��B\��<�GM<��7<!���\�i>p��8�� S)e�ʺ��x6�[��!z��׀������[_��,�����nhWԶ�Ό�v�`��yR{mԔ`OL*���=��X/k���V�P[�ħ%���������߭��\���:�:>��.�x�	�6i���e`̠�<ּ���� ��>D�4`MFk'��������Z�iY���xV�R�C�mQca2�UE�A�\��k_�0��R��B�>D����ֿ$�6'�̪9��3�<����꣙�>�(��k���>�D���k}��������N� ����Ri�˼�2
�)r�Y�x�y�>���K/n���� �*� , rR\�?,$���o&��>`3TP3�%IX���xz9h�}13��������f=Q�Z 6!!���%O�;�����>8��-`��1Z�O�,>A8��D�N���,(�գĥ�y�U!�p�kTd|Q�:��fP/����ԯ�|*+,��q��^�'�+��*���C)1�_6�Π���4���Z+#��-�on�5���3o��;U�z��t�T�h*V)�t���R�@0-6^67r�OWDQ�&��,�>$e#m���#k�f($�/��.���m�����1ä��M��B�{P0�n�3*���5K2��+��ܐ_ŌL��Pǂمh�^��;E��;O�>��? y�B:.;��P��H*��q��������^��?�O�o��}I�1 �*��H�P���Hp�<~��!����k���dց�7�'�������/P^a@7ز@��� b5��ů���%�7IӀ�(���k\�Y`�ʻ�0,k^�q�.ڦ�Cf��
��j6�4�v'�ŷ���e�k� �ܣ��Æ�}�6���!�y�`^�\�z-�cW����V�iVhl���6�Sj"m����%*���z%�-���?���H ���H�iS��,�L)�γ�]�Q����E�$��ci)-g�:K�7>���eQ +��Պ�ͳt%運���q�ꄰ=���,0g����������-'��h	C:�d��N��+��+�E�Bm�>������j�daW�L�?��y��[?x�$�������_+0<���b�9���̎ǈ�e�BzE�*�d��H���/9ow2;�k�}A���P�k�^�+��%�����4����ďqq-�w
��S_�F�����V��֕\�xc��N�r#3ɞ�11�%�����9�� 2���	?9��fE�o6��l�2��@�Q��������'|%��7D�~��P�$8X��zva7�� ]@�bƔ�Y�l��?�q�7�b�*��$�+�gJ4vW�%$����ѣ�}͏k+��<� {+P�_�I�W#�p���v-YJg8�Ũ�A{�aY���#�w\��pEF8��P�d��Ȼ�N[P����8Sf�����:��=��w���MޮR��g ��ۑ�!��E?@���nX��~�㨙x6z����}���Bd�zx��<��\��8�ȁ!!nsz�
�+�(�s�ZēԓY�J���Z|2RQ":���YY�j�.�ڂ�{�X`	�!(���IbJĆKc��k��6�Хy�m(�7�W�n��s��5ݬ�M��Q̮C� Z`��?�����rn�9#�� �$8�^9�G%lot��^,"���_!1*�˿y.zǠ�;��ӄ�HM�=va)�K�@7�}4%V��������m��	X���! z�� �N�w
0¸-�ei{Mp�&� ���p��#�.ry����}�w=[5ȩ���z΢� ���vwa\�e���?�L�XݞO�
�*�i�(`���<ܖQ9%�Ç�����>������4rյ�$=�o�U��R)+x��Xkw�,'A"��P�$itwߗ}�J�mK�!c�#I��s��D�hr�U>],�����Kg�j{���=��s�Om�
��u����İ�*�f�{	�����["8.���c��2��DZ����|��$�Rޡ���O�F����as��'>#g�N��	D�ü[���c`��؅�6g��3�& qk2+�c*��+�1��O�lZ-e�5�w/�5$���w�{�u����-]��A�0�Ț%3�XY��y���L�
?T�X<��)ʆqഛr�:�,ckr���S�O����P;��M��<N;�~�����Al�ARPH������R5�������;�M�P_s,��@�1�.H��$�)�ju|d'�̨+h�r"�;cJO�5�|�� B�cH=���C��J�c�+�h����B#���fYz��Gkz܍ݿ�`�^�@h*�Jc����`�S%��)��x��/�NP���.�%J�^QI5���h?��5ozU�)G�W����̽���Dqgˆ}��C�r��"[�Z�k������Nb]�Z��;1�6?����8h}�]�sw�ؙ��d�+9e>G�����ǃ�LhIT��?��0w��+�K�R�墇�?#�Z�`���3NK�B��]�I)O%���G�L�w�gΦ7َLt�y�t��x$��,��s}��.k�᪭{��{��rp�Vx��\�z0j���W�~�N!�[�� ���-�E^�B�&�`>�:��WT�ށ4�J��Gm�I[�ű	���R���)9̬�9�)��W}�*�u� -�3
�KB�4�~fi�)����t�q�}!�����+��� r�����E�`��c�P�O;i8�DU\&��{[�ÿ��vA�-7n�2+^��#U�:�u0�Ϋ��:E�B8� �֢�qg��{`/M�Yb�O1��ݑĻ��x^7���b�� s]��Z�糅[y������\k�I�ș�,���
;ZS����o�s�J^Zf��U����sb6��-Y�=Qd�$V4�r��x�~c�h��.y7^$�yM�����2�5V����\�[9�����_������3���MƸ�fm�t�[����XO��YXk?�b��C��i�V�A���0ℵ_Q�U�(P�_/��W��������X�0K�Ǩ��+|z�����wo�mf°��|�6wY��v�!����}S�n����V'�L��go��kA�����i
�zQ��0�r�C��h��c�8�-�|Rʎ���[�*��3�0d�܊���_��L��Z����|vǭ����أ�8��&�KK�ٱH̈́� Pz�6��NaL�@�j*G����}�OKK�I�}pP��
Ҹ����z������z�E�D�a�|\5l/�fI ���ʝ{M�'}�3	~���2[Qpr��i�.TXD=�����o�H���?[XՃǒy�]t)�@9�C��t��~c /���G>P�#b�7�2Q(i�ט�Gs2��p�h>lh�X������3�&7�$�!��+B&SX�]�̐|������8p��ʓ�/&"_��k��XO�_������D-�5���$1u�E_^V�9�I ���l�_c %�x�K��c�2�����c$��R�]_8$)$@L�.[�dad��讃b~d3�]/�{���W��5��/؁wi�k��$��$a�G��H���M�ǔ�W����MB���W�������d�g����-VN<�:��R���`d�W�8�b�WO%��R �g�_��b8���\T��5Z#x}+3�ZRϛ�
3����/B!�Ǝ�6�4f-�Qx׿UQ;��eWڏڢp=�=dy�__xH��q}�������ؙ	u�-q��Y%���>Z@�4�!�����9�%`O)/.į��嶧Q���.�|Gnj7t/��`�����s�]}C�� ��5v���I�o�����ˣW4�w@YQ�x�\jp�?�sa����F /Gdx���ă\D��'Za٭���_�#h�=<�˅��)��T��*("�f�j�C��4��r��@j�S.�̖�4�C�#X�j�b���=�G��]�+G`�.-)mS ���g�~�L��P��>r�S���3cd�չwAx�X���P�r���v1�+���m6i��z�0����<	���C��Vփ����h4&zڠ�p��N�!�֮�Oľ��X�Ф#0[�@Π��uDVǝ�M(�`�g���?2���\v��g���[�� I[9�0Vi���e�V;�C~��p���5j��ܞ�4z�yv)<?�����b���r�	q��4h���{�R� |�����E�͙��F�p�h�|S��
E��U�f�X-s�g�����]�C���{Z+ $�T���x{7izT�J�k� [7���h=�k��@��N����9�R�ۃ���9`��s ��m-K
��J,Up�pv�g��Y|/�R���>|mYdy���.@�G��<�i�����b)�^�=w�W�-�Vm�;Ia����c!�h�
�bu�����G�7��O�}�$�֫�^�`0ӆJ�V0	�(�YԴ,u�.3镫B�oL�v�P�6��"��ެ��w�VQ�������0�U5�1����m���QV�ln�2��w�GcR�LՐz�<L�[Cʠ��s�:��o���ţ����vq#����>����L q�(�AZ{�H��F"㠷�fD�j�����P�V��\R]��j5�{8H1vZ5���ϱ)ڏ6{��	U��w�:!��h9Q��r�y�o�X����5✷�R��<�M�Խ��C���]a�sZ�����olm9�HQ;w]��c�S�s&,i֮����Y �3�.�8W�@��E�ʯ����~�.-ｻ�RI�*e�ei�M��*��9蟹]/y]���'���A�fw��;�Kw��
UC���L<X���u���E
�d��݄_�ǌ��"��<&� �|�@K?![X�*�1���_gӷ@�C�ɠkf�}r�}hˬ�t�T��Fw�����
Y8]0$\�r���Y!�
А��<�t���X��u�ҕf�x�4Y��Or��tď`c�p�선���;�zX��%Ɛ!���P ���ᢿ�02c瑣�rt�~����-��jQ�K3H�Sn9�}�Tjnp��^]8靿������*6���2bH�x;+��d��h�~B��u�������sd�\:w��E{L�O��J��qf������Xt��m�$I��b��#��J% 0�ɠ���#���Hl/7��]�p:�c7] x��c�ߐ�������'�ji(	 �,��\�'�@T�Z@�ܬ��b�lq1���t��7W-h��GCs8'�w+���
�^�6VIT�K�iGhճh">l����&)�ނ���۹:Nm��u��T&m,#5��T�u�Caw�2�9��a�E�5�7푏�B�v�}�U��jW�t����q\� ���F^��ku�WTS�_{7�c\OZ�B���ɩ�vF.X�%���C���%l���|�5R<i����k�0;'͓a��l��U�O��t."�5�3���R
�Wl��5����
3�~��)��MzM��ܾ�`����z�ٌ3��I�ഴ@��@I(�t��_F����E7Jş�6����Z�)*
y��Ut�?t[��"�����@XZ��V}��.�t`��æ����_����0i�lt�*�Z���X>��^�u��w%t	�et�o�6ʙ�����`��2��d�gF�1�t<@>�;�YO���`bhv.�]9ugI9 �bY����C��v����0��(G+�͎���f2�!	���h�`��"��g{q����s����6*��#��Ǜ��S?�F�a+A��q�6l�F�7/�e�}�&*6*�K/��'3������������$?���*���!bػg�؏���3�҂!".xC:XZ�I�Za��'�h��$�O���Ū40���y�Z����@��[Yl�-m� ���,|���ؽ�)eL˾+lɹ
TX�)�1�ٯ)7��U�����:�����3����!�g���W��~�7/��S�=8ѩx�+ѷL�fS�ݣ/[9c��2u�]B��+�f�D���N ��1������������Hyx�[�XN�"�n\�������rd�޵�įP�:�KH������١���؇�à��v�� �w0q�?�n	����F�x��ՐB�	ps�[��F%J��Ҙ���l֯��d��_lIhG)�D�Y��9��X�Gy��kl�s�;�^_!=��@@U�1�jAF3j�f�ڒ���?���!�x��ZWh�/߾$-�E����?�S�\���v*W��%[�^?�����p ��ن��'z��^���#t�@Y���M�S���m����k)��]�yO5����)|�Z�5��0�/�`�0��풞t�8�Z�%�u��p� -Mo��ҧB����Ejy\������)�Ĕ(��TI�_�H�z����d}��"Q/d��)��
C��xX�E}�sظ����� o�I~:����Z����1Q��`� �㤶0�ZNބ�A\~G{����� i��2�'s�W.�r��g^�#t$���������h�3v�Xe�q����<2'>��+� IYj��ͤ.)���R��&y�j��H�C\��0AB�86O���Q���Jװ�4�ҟ������[!p<Z��j�N��߽�`�gP����m�̊�]�l)�Ҕ��o��S/YU��7�vm�h��c��Q$^�&M�������w)���=��j��;���!�!+�$����︢ʟ.�
I��r(h� SӴQl'S�)p�r/	Fr�a7n?�V0�pۤ���*�na���Kl�� 0D��
n̎	Y@�����d���ʙ2�������
�_�>	ĝ]Aq#R�w�M֦��v����#N��X�Smk3���E��>�ʀM��i^���kd�����f��J����-w,S�k
�v'�$i�� E�O���8�wɑ՞a��a�=�o)���C��L#��w�~,j ���-��9�}�S3��ڛ"׭t9P-1���}ǣ0���%h_�m)��4��1⇪��g�NX��;߷&�̟-p���8�+9��h�������˽�WfR�=/;�Rx�M��#JQ���-�o�zG���NZ���1B����Ӊ�^�z[����"Ѣ�wWr&���k>���P����jj�H�V�F/���~U3�����,Qz��L��Z�
�K���ڄ?�`��4�b=qd����]2��A�$���/���L�ˍ���,j���H�~��]*L�����Ӂ�������/�9YE2`g���*\9�xg'�D�
�r`Mɐ��i�����?�ߗ�3�m>5��|��ܥ|A�j��P!#`k��B�G%��w�(�.շM*EH�'_ͺ<�p��5k���6�n�-v����SE_9��R�*�:�h4��]X���*ȼ��((c�8���,E�AG]�ݗ%�l��ћ�Rl���R��}�<� S��g��wLxI�]	j���)yh�	�8���^�*:�@i�8ğd�]�P���aʔfd�<	+�r�OLo�c��Xu��w(�^�	F�~VKu�u5E��]u�xy�q2Xz��`�ni_����Y��`��r��I ������4�\���wͻ�$�}�I�R�<���{�Y߰[��,~�w�t�U�=bb<ls]�ע]�����0�e��q��K����Xk�i���2�������3�N�����1��	��!��)IM��� 5\Vˮ �m�`����>��=��?���A�3|F����!��/�� u}@�Ǳ�7����'W֕�Z�?���J=\��[d���X�N
��{�J2�Gg���3�>A����+Ĩ}iA{m��8�96���0�7�(����a6u3/��c�>���Sڳ&B��_��e�G�H�/����X�k�(P1�� ����*?��4���f̩P���[��3�s���=�z�ķ.D�6HB����x���)�	&����a�a�Z�=G{S�2�7B.	��I<�X��y^�n�1��2!ά%�wj��F�2�.Q&�5=�<��o�K@W�ºc�m�Nw���1�QD�~���X���0넙/{-fm��Fkҟ�w.ժ�w��,���Y0�ˍ�]���CR <#�92��[e���;�&Ю���w���V� �C|����>ެ�晗Q����S�u�t�������|.��A�lD�#������H���'3e���!�-Ky-�5q��޽�F���#[�R����'�gE.J�X}>>��#X��֚ѳ�J��Mz�)|���
bb���}���4}'MG9L��+�}$ޜ�����ݕ��P\H�Sʨ���;7G�m����t����*Ϭ��/"�/�T��Ȧ%���s
�d'D�66Y�\�ͅt��EX�:�V�>�"�z�+�]���ǯVlm.tL�R�J�+��Mog�������J
�^�Gpe��$L$Q�1@���kL�w���b�6���#y%ń�N��8���6��q�T|���8��[{��"h�u��,�����"���)��m� ��OX��:*]��Z1n:�g���v�w��Q�-a�\�!���[B���#��*k�|�;�
Һ`������n�����tg��+�͌���ؗ����L:�|�>�r�Ϳ����G���%t�x�<��۾�����`Y��BG�yȔd�7}�u�+AC��ȕ��ӛ"OAZ}!a]�B��I�������J�� �im���8�'	��@D=�2������Bi�����X[��̴d�͂���L=��X'ڹZ�)�6(Tȟj��ٹ���@@�N����p���[Zs�%@O�9��Ϯ�2��MO��e�n�^�^��~|(��tҒ�'-���^1�f��$��e��^�k�9���f��W�P3{Qx&��.�Z�� ��6Vr���]@Z�yC<.�{�'zy�쫅�ݥ����>�uߎ��#�^�z��in~�D��;t|��_Σ�����yMb���m�4/���qų�t W�u�<�u;ø�W=s_�z<�Tn�媩7i2��n�B�5v�>H-��� PW�u S:��;� I��,v)D@Z)kr#2΀{�+d��^r��l3���*y3SƲ�x�ΐt��C��ɅrZ�X�Oa��T5E�䣼mJ���g�-�E ӕ�w�51(�_��� �،�}n���i�(�xwn끷(�+�|����D�X��]
J{���-/󟎌B_�]l�d��A�&25�sՖ\�B�,
���	���Z�G�5��*��^жho�����#��Uھ�4ᧃ���D�x�P��Ў�(8F_:q�fXi���O�wB�q�Ynစ�O3�-�]�ҵ�|!�-8���L4�u�bH
 �e*��C��T|�ִ����V�pJ�n�r�~;��0�@�5
ҽ\�L�Q�'�S	��If�V]� u���*�)yv5&V佴d>����;F����z��?A;+���Ҙ>�#��E��a���;�#T�%G��Ab����u8��ȋW�쩑�Z�"����rJ�R��5 �$�����v�h�'x�Z�es���.-��[W'����~�T✧L��M�h��sޑB?l��*�����D�v�
	�1F'�\if �_��|m܉{�WvFY!=�'��$O�D�}t3_Ν��t$��#H���ct��2�iৣ���k(L�̩��2�k����73^H ��HG2�fT�+�����)N8_o��Y�����J���L�/�A���*�?��Y�k8L����~a��pIA�l̊6�ή��4;���Oj&@�Lە�yS��)�Ip�:ɴ��)�Rs�^��Ͼ�P#hd�l�)}��p�ڧ4wF+�نeӘ��2x���E�R�t��BzQ7��	�/4�&��K��!�]�g�wkJ�,mͬ���[��aW/�w����o��v�sl.��E��_�3��[x?D����R�ā�5=��s?����;!�_	x�EW�c[�9!c1���r�G�����Uqa��{JS�T�pђ�Vm�)���<��_l��ƻ�p�B���H��-V�5,\���~�x ��OX��Ic`�75ty9�D��!.��(���J�z�xm?�|��<P��ñ%�U��� &=tX@nTi��*9�p�7�;%�	�L���1y�8x_W\���O��Q���d3�@0�}B��b�K�Zu�4�w@N�ƃ��`G��A��^���i�A�4"���s��?�b��D�S������QRr����i��7K�1b���$���`��7n��3���[u�h=\�j
���BY�("XSF���g�q!���J�^��6m1��T�m��-G���nJ�~?A�[����6�n��u>�4����O&��ϫU1�ډ�5�=�F�ş�+��!SoH��������y�B	������%�[]�ʃ���x���>	o��;�p���-�JyUQ�$:΀k�	���0��fZ��B[=����.��T�H<Π5ҳ[k5	5^�,�I�S���e�q�-��
<�׽�*�H}�?�G{��캩��hw!�P�N����Q�"Q��G�z���J����T(��j����Ձ�[�u6q�-�	��7������xl�N҄+ꌛ�/'�?]R&�(���"�gA�-Hw9��9<��#���S�d�m���:���h\^�r��Sh'.�U@�F4K)pP��n)�Sۘ&��U_t*�:d�KO���q]���V�׮z�e��G��f��k�2ѿi��B�]�wAIpyFK��$BF�zνC0�ޠM'ł�dIq�#���m#�ه��?n��F����h�����Ni����^��5�æ��~k�`�{��6 <�D�fY����f�v0�j/���0�J)�'���d�i�f��g`u~����UVv{G6"�dB���Tn4��r���x�R�? ϟx��ī8V�����&���a0�`�"Ȕ&K��D �� ������5�.��u��qJ��¦��Lycjo�O���9�[�ڡ(��6�e�T(-"��!�lu:"l;�o���*o�6�,�C�A`��J�4콦�p�����b��M���i�6	Li#�Czb{M@?�|*���P�:"S{NL�U�b�Q��E�}��M�Dժ�ܬ淅9�_����V0Ȅ����I* �	��tH�'he
uE;��n� �z	�jҳ��C��#�	"$]��l�6�R�׮D��X�С������$t[�y�����zQGNm�&��;*�_�,�1�ޘ�+ĭ��x�(2�е�P���c��7�����$�/}�x�P
p�����Ǒ9)O���h�	n����4�Q#�j��hI��0V����(O1~ݕ�.����sW�ģKV��c���A�F!��L�$t+B���"��׏��@��=���ҭ�r�~5m�[�}Z��C�h�s.|׸�Y�d%n0��u$	�$"��ȹ�n�.���Ae{��A�@_4�3]�|͈q�%8�<�CkJܹᚋ�ޏ��4�d�UY�x���ؔ�狙�S�������d	�[6��	���p���Lu<kQ�pL�maP�(�_�Ͱ�����ż�&0W�ԍh��M@�ί�_�˺��'fV�f��b�E&��<��G��64�DI0( �lP< -,p�G"�	�;[�9�}|ﶠey��S��i�x��}�f���`Pmj*����j�H�O�jL�_��yV�����~��\�4J(BKB�=2R�I�ݓ��-�B�48���v�k���(��-��"��$�?{mv*�v-}�ѽ޻�nm)�ʐL���D�גWgC3S ���mSU��9PX��"yG>L;��������/j :�|�6����R��^��`*%��Q�"G�-�_X_�I��.z�ݫCk���˛�6R��r��0�T�@����qF����֓�77h@��$%�nL�O�;2� ��+�]����P�6�x!�6:�� �h��5i��S�������.n�ԇ��T3���x�����^�o�&�KԴs[
��tQli�Jl-�Am�F�Q�2�n�#�Z�JWAY ��XPS��k�F�{�
9�ݡ 6�I,B��Z��{������@�d%�a!�Д:-����f����P���z��W���6� �x�X��g�X1�/���n<�Z��S<��b�*�Ͱ�ow�w�
x�q2[��~��t�39y���"  �F!A��5�� C�H�e�hz�I�f����׳Y�2�W�������
�����"+��9�`/7��#������RZ8�g�?�!3�*Oӭi<?G����\+v5N�f�e�Ȍ�-͛f���p���3� n�@pݜbJ���kb�8l�X`��ޠx��݄��{]T�׈�U��,��o��f����N�Iv�`M����Ms������,����ϕ���xǓ�Q�ʂ��8���yˮMY��7��1�*l5_����لȠ��J�������� m �Ik��x�&r�tcbu�hp��U(�@�
^7g�*�߅U�u�o�ߋj���@��jQ���2���D���L��w�hŮ����ֺ&.S#WWxk���1����/�BY�
'�{�}3��.�!Q��е"aIS����2!��1W�'����(Ti�	���u�nfg��9�)�#dߍq�(��F���3�qptm�{pt;+옙��_u£�'�sq�;I�f����\Ro�S�y��į[��
:�T�#A��<�щ������;��*��}{��?qd�m�q(��W���J�v2��9|Ѕ�l�a��0� ������Aܺ�m�xή+NY��t��©�Y�L�N�?���0?,�A[�=%rP!�P�w{�*H�r���)�x��"f�G�nO)�bfP��&ߞ�k���B=qa.��
�}0������iYT�;�*D�����4��J���ӥ��9*����W�@%�_&$1&������h.u�qES��xN3��~ �Z�>bu���B�}�='���b�%|T�&�������F^e���;٫O���Kf������aFW���_Q{�V��.QW� M�^m�w����W��P�S@7U�$W�;���3�.�A�X|2���<�ġ/�Yt��l7`�߯���7wu�(6�Ey	�t.�:U�K'V��]�At�2d��%�N}Ch�g�(#y��i��l��/���<��\������� �ݼoBˏ�=�
�����a��Ca"�K]�.�� �A�H�:�� �aE�����[R�NL���X�J؎z�_�i|�v�1��O߶)���n�9	P���g;��N������+頪��|}}*i�b�$���߾��K�2���=��g~/�2�&�����d�+Q��8z�}���ݷ��R���5��!����A]nħ�O��s	�Y�T�L�m!�G�e�{pL��e���/��m��eՓ��v49�1�ތ�v2��R��,��0��{t}Q��$�dml���D���䢜m��y��+�GQ��n������"��a�?��e=�Yh8��j�h"R�q�����6a��_vTf�<���Q��[J2:�ȿ?(:`HiШS��jNl N$��''+r��r|E���2����t��x-�i�����cy�x' <<���.*n^c)Oq��O�j�4�N��㡃pl_�����Fc��7R���2�g\~�fΦG<JzU�-����uǣ����݇[S�9�u�xN�V
uF{:�Wi.1lDQ�����x�"�1�oj�!/��Z�mz:Tn'��T��z �:tׂQ'$�����ɩf�@{��x�p)n##�z1����H���7�a��.֔X��琙_o��\��v���{n��t�&0B4�<`���k��������:�@���˅*!�k}�k��{�ߣr*ڪ�'Cd��W��z�Q'�+�f��U�ּ��St9U�+7���k�&� K[��iƔ.��ҝ$K�8�]C�k�k].������px�?�|4�M���E\��Rʮ�J���w-fM�Y,Ĕ���Ke��,D@�4�ָw
�FN|���-s�� �6`�>���+���7��ۂS}����w�f�Ci�}��f,`ᔾ1�ǿj�r��3`M�����"���آ�7,S����<YA��w?[b���mpé
��d�����A�Ib��;s���8w3��F��"�r�tb\����h�DP�Tv$5��i
z�($A���3pr�dJ�oF�@�X���/>?�Fu���Y����3]�������6�kp̬�|w3��Hi-i���K2~��a4�f���TT4�P��=����	;�x�w��Y�p��t�:���C��
��V{���F[Of�\��>�tc�'�y�wp��6�	�7� ٹE/[c����>�e}+]�W�S�1 �!c\�!b9D�m�3K�Ҳ�De5�nR���Sax�~y������A:�S���U����A�+�+��0�Y��&)���� ��m��8BX�`~�̈́@gE��и�D�_쥵�����Y=.���zX�Z~
"�퐟�����<e\��oU��+|�\)����M����c��F��]=:�d*�t��d' *�Q=���� �U�Ɨ�А	�l��1���SD�އ�eֹ��A�5.��M�6S���U���������ϑn�r!Ș*�BQ���j�Z!�s�x�LGDO`W���lE��:,���^Ą@)��)��K[����&�
\�����J��l�j%Z�Cy�Q�~���N�M�(�n�A�$<�Rל�H�ňW]��&��x��_��'�iϯ�+�Ə�<~y�c���!J"E�k�P�*���3 ݢW
Y���X����|�ͫ���U��㞁�U@�XL _��8�o����9u�������&G��TJO�	�-}1�ޮ𭐠I��0��pB�e����G�yH����~R����/t���-�٠ͧuڹ�	�݂45KX�DŹ_El�au���s��,�X?�G\(�#Eه���n{F�9x?W��\ ��5�j���>������j��z���罨�L�u ;���j?���3%���Xpa:\	�}nl�R\u^�&�~17�ظ�O����蠱V��~��u|{��ݾ�g(?T�P\Eߗ���ϩXU<�)�o��h�R����e��b����\��?��h�{/�#�Z(d���n9��~�����{?k�K�M�lᾜ�]��PZ�vj�
�%��h�V;����o��1�Y!��VבoSMw�����<I�K$��L:�E 
��U��1锜��S�+�td����]%8N�?�م}��
��G���[�n�
r�|����[�_	�Pc��4i�+	�����{�K@-@7�m*s7�,ޡ�3X���p��YPS����2���5�5P�2�+��ݗN�,�A�򲃸��� �*S�����p���F�`5<Ҭ����p���f��ݝ��Mv����g�C������֪�1H&9���0E?�j&�a|J��'^+���
����*m����ޯ�}b��qԮw0��~�q�6� 8����\�M�޷B��Oh�LsfK��\y뽲A��d�ɏo�8���+]��s����AB��o�8��EE���p`G� �!B��x������@58�d����%`�EDs��=a���p˞{c$�Rq�||�XB��]���2�bh�Ax����W��S]+�i�G�eZHe{�2���� �$UPI2HeG#;��م@�i���Y=8��ހO�0'xy	vd�/ZϲAv�P���w�\Enߔ��C�����m^K
9=v�~�����zm��Zh��ۄD݄6���C�qCX��^H�hv����S�B�]�P��Ii^���͔C�<�<��rz�*�B�S>��܈�����$��E�RW�4�+�{<Iy`i^����v�;��Yp�Q��[8�	�ȑ�jd���P�6�:<N[��O�!q*�M ZG/�{#�aI�ڠ�?�8����=a�zw-�-r�Ʃ@���(8�ߋ��,@�����'����w������D��C�E�ǈf���0S�6����%�T�X�ˍ���`��ޫ
z>�o2����8ˁZ5�-���q�l��9K��΍���w���TӶ��J�΋����"憆K�͓���@�p�>��'���m��d���a;��;�G}!��3��f�n|1��8[�VW҃ZY7HWPl��&��C-���`A�!�)�WV�|r�_F���XF? �F{v9RB��Vw/��_�f�Ǉh�-��hĉy؉$sS9��pԩ����!%L�g8 u�'��;�̕��kl���)�֓�Y���Wh~0�2����bЇJ��Ò�cj���A�9�`/���A����kR����Xs����$��?�|c^�����R��:̓�:�j/�۰�a��@X��7����@���y��b���Rj�B��P�Ga��J#�n�E�M��h�}�9{�>��H� �S�֓��,�*��̶% �5�U4@�%� ��a�:^��:0PZly�9l
5ً�s���@e���y���X��:��W�1lz��E��BЭG��f~eD��xh�ܖu���#�Le&����:.qX��>6о����tRi8LRŝuG��Y�,P������U.��~��h]��{
�fU�W�DmTbvrH-�#A ]�0��x���$�B��8�U�ЂV�B&���D���1�e�9G��-c!`R�$d~x�Zb�^S��/�3�Θg]W����Eq�����^Ƽ�O���=x�U`=쉳#����8��d���<�d���	��?gd�6@��O���V̘�ol�zE"*H���60}�i�^�H�3�����(F�#�C ����?/�%��/���=�!"�T��Nj~F�m����*�����S�ߘ
r;Ѯ2� �W�L5EvgW��rK��=�WE�����]ܨ72�"f9g۳Nw�:�w�u�䩈N����A��Be�*�p[r��:d�e>5�\ÿ�X���8|��+�(��kE�xb1W���1j�<�?6���R���<n�Nռ�e:Q��i��bT�l�Z��|�{lD�w�r�^�Y��v�Yґ��޲��^����6~�]��$��ho�kd�36չM�\X�	g����,�sT��m
���	���5�,�qbJ�׉���}�0��;�W~��8'�b�]D����cP ��ʏ����l�w�u�ym�7Қ#�%(MbC��c�Jh������6��;�8j饠��J<=/��|d���	V�@͕�,~ �C��E���U�ז�rl��O�$���2�=���-a��3*����љ�����b����q��nh�(�������	5\�v��֘.�KݠÇZ_s<z��y�2H&H��DO8�+�}CrR�&j�Z߸{<�_�^_�Y:my�ei�
>�C�ғP��ؖx�JKc��'>B�D,jc
W
�.dn.6K2y�n5jޮ,�w~�O��p��[�����̉87���å��f�!��\~�"��ǔ�9�+	{�o�A%_����>�����SD����e�(�EWswR�MF0���q�YSb�[�+��:qO��9cZ��ӯ�mI�%�����0E[�� ��_>k>=cf'��@5X(t����^[�>y,.��<��5�ׄ��_������$�.�qU���	��vd��Xe�����!m�\b��a��~�T`Ǒ:� k��o�rM�Z�z�1�X�Ζx��%F%ǅ��Kގ�
` ����9f�=d��u�ٶ���x�Da��ۚɱ~).c�� <��߷��>��ǤFC����+�z��eE{��c�X�܂۵'7h4W���}�@���p�D�k�!>��#�Y��	���QnM�hוt�B��f����k�g;:�1]J��D�D�Cʁ3�Q`V�CY���5���Gs!q����eV���τL����?�r��D�
�#����C#E�d&���x���=�˂U�X)��<�n��G]b������ڏ�z���
a�<W��3�kܢc�K+�A�k������4��O���`�X_��$�Eqtd�&*�[��U|s�շT�l	�|�s��k&���㲊�b^݁��2!T$�	�N��>���3��������
6�;��Cg4��ܔ�atq�6�Q��i����5E��Vv�+���Y���D��V^���(�_�Ý���W�-Y�����Q����^iټ#>�(���W���>��@K�R b�.�R������-<u�,��j��L��ʊ���G�Gы:�OfI����(XdX��J0�o���y'*�k!:0�l��bp�����
s��/;�rn0s̼���	����P2X��3����Y�`��"������8(�[�R��!�ɮM%���6��Π� �l�*0.*u�9�c�=��{�����e��$�mz�= [�T���i癗�������V1�����q������E��qq�N6|eZO���J��~���J��<��W,7Ӌ��@bk!�ح┤��㊴�dr�N�U]{z��}{�����3�aSC6d
o�:����A���5�χM�J���f�&*e�b@��;��J��8��vP!Xd5nc����+&`+���I�ưeE4���m�D+&0K1ҍá��y��o���%�Yn?�JO,3��%���]���0*��JP!lCؽ/ȃ�NoSVMgg���� �� ���6��J;�qT��֚2��Յ�u���h@*�HY�{�J-�F�m�BWKV��s�V�@R.���\��;8��v�~�]�+7)ā��AjM ������\~Pu�Ϩ�o���� �ޢ�a�'9�$�7��5ɀ8<�#���eu��Z�Y�0��#n�~z�	8��.%m���@���%0t^DzQ�/�� ��8v2�l�;�G:I&��j���}�<�m-7P�5� �x�x�������0H�L�p��������AYC���ސ y�[�c�y���8����ޭ�8N!H�?� (��]���>VB� ����,p��5�?v����g�~�"�ߓ�u|��:*@v��a���5���Rե\�q@�8R}�jNv�a�d*?���uuu� ��e�.�o8��[BB�Z�'͟��n��Z|���H�OZ�؈���f�b j��a�G>p�ⶽ��d���T6��j)F�U�H 1
���L8 =�.�h-��y�piT˾����+8�A��J7tq
ݺ�o��]�~,��πc
j�0!M�D8�1���%bt���!o��T�7�>� �u�`�,�t=���f{�B�@�ԠGּ��c����b{�0/���.�Ke4�\��jս'v,g;R��֣-��
K��L>�Z�"�%��W��Ô�A��Ƹ�I���	�S_��F���jt��R�W'��!`� �u�?�����#�lU:{&8M�ү�����/t@H�2����J{)�
\~�������+�����7�c!��X���P��>x^}�M:��r�~�3�Y��.�Y8�h1����O�����f4�!���M�9�`K^�i�x8k��� �l�C(��W"�ަ�x��)��aQ���P�"�{���V�`XC��4s�<�\n%���=�B�����ŷ[�R,���*�gb��6�
^z�Ja0%��]Zs��/�^5
E��a���Ќs�K�ZN�r�o�*�7!���Ԡ'�PG����&ˡ]�A�}�x�����S���G<��'6n�*N�U���Zc�>V�
zJ�X:̆�s�j���2�!+n쪨�k�n�~� ��p�,����%�Ŧ�03��.xo�%�;�I˶�v� 'P�ֆ7�冞}c�ˣN~��f�"�( W9�����M�~��;s�;�(nL%�@��� �,������?:����m*���hrx�(����Ĵ�_��܌�4���p;#6/Y�*em�	�H�,}*��zG�����=�����<�)�*�X8^�YZʖ�P��J�V�S�̀s5V	[�7�X��AJ� 2�<��|�(>n�}eFy,6�	J+�jށ��T��"�31�`P�bߗu\��x����E@Fq������w	B��2$?��g�)�8c��x�����^�;J� �8������U�Qʃ�}�,"��B��oŢ"�|J�c��y'Z���H���'���� l��f0��F�7ث@I�\�g4GP��ޜ �NݰE_��կT6�N0­���5im�Q�<b��G�8����z�=� ���X���ȗ�8��D��`�.�����|m	�:�ΑO���W������7��B	q׼1�8��9�"o��xzF��`)?`в���krE�J��-����PVE�K���TB�ӝ�e����ؾT��y��(�$G����U��١h�ET���[�ɨ='O�ov�����=�+E���
*ͯe�X�k[h8n�W���z3ӭr+;�c����(���h�k����$3�Yv�!�La�U��H�
�5&��}�|��Ɏ����u���>^�Ӓ>�8~�-�������oҬ��&(��%$�>:o2>���i6S�Z� v��%*��v�g�e�)GS%�O�ss�ގ�Mt�.
��*tz��l��d�9:[��͡�>�j2�MO,���h�mo�B@��g`y�m<W� _��X�4��Y=x�ǧwW�pS�h�πAdw���8��k�G�)�م����2E���C�xE]�A�RF�6��/�Gj��c��r���I�#6d�
;���"�d@f*��`��k�?۶`N%��&р������>3�+.N�^h�#rF�h1�Uu�2}U�l�Ƽ�ʭ�@��V�u�T%+]�85��蛨�nz���	n��8~�[�+�LAI\�n��5�z�z!|�)	�@���9��{��A_��y��J��}Sj�Ǯ�����h��G�U��.��<�,i�#! ����h#i8*��Dj8=�����s�EJ�詣|S^DQ��)�ñ���	I^�k�!u���"�P�Vez�f�-t�M�El�����R��솖��K�0�yKmU���ۥ�v���dߤ�*��Q4���^l�㶋�U>KCr��泲�kPD����+.r5�T�~��N�_v[�|�%D���l�0��6G�H�_���e���<�3��� W�<R���̔7�����m�
],�M�ۑ9�Q���KSY������6@:;pݙ�(�;Ǖ�Kc���]���ѝ�s=p�(E'�L?��E����i�����"m��D t˰���&�!а�2p_��_lx�yg<�v@=�A�Y2"(�VLB)=Q��%�m(���_0�
9^^�I}��))�+N���`P��_���� ��(q���K���Ǿ�S����n~R���zFK�ST$:���}.�jB9��,�$�լ�X�ڌSf#j�e+vB`b��Dt��srTwS��g�D�B��z��Ù��i�;:oY
�h���׿�އ��"��}��'yʅ����]�G���&� �D���"v������A�S�X�dΥ�j�8%IuSX:�O��u�����]�e�4������)�i7 ��&9y��Juz���e�%�.AI��e�OB��H����l�杝>�8������h�8�=K5���F�����- ����J����ڋ�k����~��X����)yt��j�s�-�}/��Ǐ&��+���_K��(��"�MҐ�5=�z�L@�`kq����9�.�<)�B�q�Ma�=V{sԶ���B�-ڊ(l^IP�:)+��%��� ���Hܕ1ߺ9bJ�#U�v��/��5�D�k����$�+\pD/N�3�4��%�oZ�+8��`򦦊{�q�s*&qN��ӳFf}���5$%'D*�׈qao��H�`c;52��/I9 &�{�)����rC�wQ�w"VA�潒��&B��'ŹB�W����v+�%#[���ÝXeh[��]�5����R\���V>�������m)�i�*<��$oY+����VI�B��-~���pDTl�Ǐ���n�8����{��+�����/r:�\� �[�������}�������))6��(,n�Y�-+��+Z�m�Xܶ�1�N��{��k�Lk�P}T.�s��"О2C���T�*/�nl?|bn~t��=Z#����,�l���E�pU� ݇ƪ��ُO~��NWF����(�s�	B�ƚ,�~g�{Yg�$X��f�]�as=��˩(@���W?#wO����]�M�(dY2��e�h����K�W��x��f^����dX�l\�_�Y9uI��)�^��qs�+H.�ێL�O9V�Yq)Q��Sv�#���ˍ�{�
��2��+?��ix1���,/��z�)���|�Ws0���;�g5��RԿ�?�-�Q
s��#BD����_Y̕�+�^P���Sm���@��=d`?Ь�U�0*b䶔�����.p��pƽ4O�a��ENNJ�g(wgd�>��b�X��ش�.�k�b�~����;��1��~>\�M�c�x�,��T�W�F=/6���"����@��ȧ��L`oM�XS��z�������7l܀��y�u{���,��`|����Ȅ��g5*���p��'.��o:ix���?�b����8h���>���C��C��?l� �� �Pٽ%v�L|:��Yq{:������f�d;�O�.0ʆ-¡hyҊ���7����=�|#�[i3�S0I .�VK���?��8��/ߊAx.�E]�F��SA��{�h�Q����L��/"wsp`�؃�_����J%y ;r�/�ޱ���Ϝ0��C2W��RM;�gp�7 ���3�����2�~��R����Ql��-���^���f9a �"i���ֱ�?X�XɜJB���T�u�m��1��!bz����@3��^0+.�jhe�s�RZr�m��	����Ő�[��X ������؄��(����J�$�q�,l��y����&L&�ޘ����j��s�D�[L�p���[y;Mh	?vH>`�/�\}���y\U��8%�z@6����G�[0�1~r��w9��=����3��"�?������r�_�0��D��uu�k��#s.�h�˘�L�C���ih<Cds|�Z4�4�P.{d�%��w���E6e�La�	y���V-9�	\1����m�MQ��""K�Y
�H	0����$jg��?�#J]]���%�A����~^ln�)@q-� �T`��&T�`�l��wo;���� �������L+�Ǯctszv똍|v<��ǄL*�� �w�M�	x&M�;���t���A�v�G
��Hz�3��|8�π���b��іc(u,7�z�L��k'�"��ݲb�Y~�KxMg"�
�M�6=ܮ�X�w�Ŭ���]7I���[�dK�.�T��lӯ1Z����G�]*�p����u	|h�o�&ųy"�H����mS�i�n[ͺR��&c�a��&��ܶy@b��+��.IRJ��'1:���J��A��j�Od���N3�I(c��aď��ȫ���
N6yatLS��Zn��՟�z���K��m��knp�k]�t��[�g�&b�Y�H�y\�#�>3�o��ҽ�@�#h$�:N�;,p7�FOn�����9�V����8��HOE�L� !� �L��l�C=j����z6�f����O�HRB¦K�m�$����F?��M����1�;�� N_?|���OZBݑ�Y웘\Yn�:A��R���F�-�	�}+i707�EG͛�2w���\ ���}��@_ic_�l�n��[�+�7�V�CY�������3} �rV�?J�U}K�����A��	i��q�����q\j��8:��B˨q��'z$!�*���q��u���T���VK�{^^���c�)�����/�	#�k�#=��&djlM�4<1I�Ka�K�z�B����D˟���t���Ked+������wg95�FE�$.�h�Y�.�BH%�'$�?��_��iF[1E�b�#��>��DGI����m�p�.��^߯s�X��\LTАd�)B`Z`Sj�&�^t��EืA������N�(�Ԑ�φ���<���h,����.��̜\��X���3�<y�J	���=���:t B�¼i�Y�P'�13yR���IO�1⛖G�)'<�ޟ�kK-7�,�d[$��*
R7�0G���V:�v��ަ��>�eX�Z2�������!������)�*�j�M�޵p:���,�Է�[N|f�5~���dS�W'��?6�ቍ]j���Vx�K|	� z��ydУ3��N��au��Y�Gh�3�����:P�����	/+ˈô�>#��<���w��L�֨ϱ�uj��G�p^A�ƑI%�N��H1�h�Hq2��1[���+��m�o�鏿l����|�/�5����
/U�q:k9�vZ_;
L�|�������^9��Ԡ��5�����L�7q�����#s�'�D�{ B����(!!���iG<�g�w��W[Y�;cc̺�Z�H*������=��ʉ��z(�C1MMyX�����PqQ�d��o2��񂟋h����|�Bj��`�F�������ݖ��[h�S��[�n=�����])!DXϵ��5��ڍb�J��+�1g���3$�p��@�G)#{����N�6*1уh��Fzem0I�2�����G�C8ˊN�����r��~�!^\��+�D���Rm��t�1��ٮ�}��jq�֡�6�lޔ,)k}Gh����w�,X�^�=�����\SяQԾ}�G��L���X�eC��*��.mwR #k�4����V�h+Dǣ[۳�u����:��a��Qع��"�{;A@m�����(�袲w�qm|y�8�|�F~*�qP������QtPu��k���G
u��4F\}a�J�*;����ؾ��m�P��yw������Z��8i�HݧHG�Y�'N�g*D��p�w�dg�K������S�6,4�*�OơX޴���?!�'Ry�t ����"r����T�����"r��?����K7P�zM�<~.�����D;����I��P9B���5����0Y�����4�)�%hP>U �t�E��`�hm*��o��g��{�iٕ�/ݝz��ʳ/��R�����G�48��؟���7���0<*^َlU?�|�Z�����e֓Y�O��}��?�Jl2�"�����*͊�ф0M��z,��H/k��X(��������x��).����>�#����Te��ܡ�ڔ}k��r2�q~]�s�};@����7�CTI��������E��?P3��4X�#�-��gg�׭�l��L�mND���l@����~(zw��x��L���80�6�ͼ���cVAS�g�4ʁ�'��?$޼�gV��'�ؾ�s��<ih��/���_ʬ��PV�I���I��{�8��z�#�$>ed���;s���� ��V�K~V��Qm�0�c����D���A��^L��6��0?�[���/(��.y߷��o�n���;�/w~�|%��dm���V���/|����ÂD�a+%��{i��ͶV'�q��p���ǚ�ˮ��5�5rL�_��[b;�u�:�L4 Ƹu��M�[��X�/����Έy ����l��B���"��JC�W��G��ɻ���)K9,H�����f��[���uH��Y����2��2;:��E���.g���NS�C���3��֐Ź)(1�&1���C+SK����v��_	��Zd x'�m�m���2ZT?/��x���y���	��h��i���"��9��8n*���':��dH�1�TXk�^����Qa�".8���*!uf�r��נ[���X��q�(-����׾͸
��m��[���s��֛s�^Y�28�Sa�	@-�'Z~i:WК:�qIa.���8Xdf�M
����+]W>hj(t�R�������Z��S�5��f��K8T�bg�W�%�F ]����\�n�Ъ���[��b2*�w&�׷%hkP;1kQ���M��%_q 5yus9Â�y�)Lޜ6��\��� t&��D	Y֊�dL�~KfV��O&��� oծ1�r���d>&R�T�@Xs�E�`�����l��;O"~�T�7ě*�=!����.�Ϝk �ñƦ;������8�#]�s$�n���݄�צ��Vw<���uc�/�m����u0�4�O
`�d*�G��
��8�-txSI�� UɊ'��+��݇rt-	UZ�S%���`�h���5�%��t=nΫ$�heUՏy/�g�C����#�C�Ax�m,2�>'��}6����Ħ��:�K�7��1��Ӕ�bg�<Jc��K.[�8&�`X%]M����y���u�"�e�O�ޢ,�q��2�� �]d����LO"���^GW�%���!^(>�����k�x,�._h�`XP���Y�~�Z��j�k�N�{�xՀ�x=#V�2���>/���m�Q�X,�Ed$i%�CtS�@?
-Mp.����U�/��{��: �>1��U
-
����#z9@����Pj!�O�T@�Z�z	�^xSx9O2s6ׯM�bφ��$9��p�^���Mo��8�C�^AQ�3Rrr��Bz;�m��\�R3�ۦ(:*�3�1�^s��sM߂G��wI��w�j�	���M���te�C�u�����W�X�]�K��
6^Ѧ�Gφ����o��4W���w�5��G�W;�FN�Y�Z�{��u*��F\����j�
���J��;S�6M)����r�=�M�� >A�E�g�}����p���c�l�2�ך	���];!��շő��O�5p-��ų���U��P���ܿ^7�ACw��:@14"�����]qEդ�s�1���W6��&�L߉��%j�p -�:�t�VL3�5�����6ѧ���k��+`/����P%W<��T�H�Q1VK�b�� �����-��D�F��كbɀ�_E�s�"��@7�;I��=D��S���B�(�GA2P4y��Tbj9�*�K
s�WMƆ�H<�U�I��gbm�Ë�2_�fd8��K�R���7����
����h�����4]�M���0�����'�U ���Y50�e�Ր�I+��KWUZp7��Ѵ��8�k�i�S���h���)��폁�s���c1v�(- yq�A����q4�+i;x6�4���"��Q�W.<^X�Y�`F��NG��5�CK�:V�-[�5�IZNQ�icŕQ���F�`��
h6�[KȜ�?�ʋ�9�uW���Y}�;���VV�~aI�W�;O*S(*�Z�&B��7ڂ>�4�w���%;E��w.����²�py}:�?�I��{qv=��_��gXSK����J�yj~L�m�:e5 �?lj���&�b_�<@��ǯt�l�gy&�zޣ�[�Q�Pr��<z���iG���4�ty3UY��ۍ��X���nu�U��Y�q�������	t�! [N���JӜ�6�TT3�YVTT
��Dd�I�$�}*���T���>�>Tb/P�@���eQ*G�޵v��O��c�u1��YG��b?+��9��9���u�g���G���z� ��H»F�NZnkǣl��������t
m�l�:-T:�4В��2��������KJ����\{+��6�h$7o��ׁ^�/O#f��t�A��L��
<�*n�:�;Lת'p3(����Ҥ'٫��Q��׫�4 ��L��q�4���囶��&�1<�2v��ꃻt�}]����C¾���e���uNіV�*���	�u��g) ;���݂�C�(����NOpuM�[e��PWSb����%��ެ�\�� �20?���0#m?4|YBf }c�V�T-�����)��6bA��^��	�Lx�tƝ�	���>Z�ꖫ�Q� �7�R�ahZ;P�jӞˮaXUEj�rV6�A;�Q}�����\K+H�}���j�G{������ICF������Z�����7�<�C�̣�%7]�d[��,Ay��L��h���T��d�@�3ڋKe�4�:B���2���/wmb���m���o�B�O�����jVR[8�d�U@�7@�ܨ�l�6����E0�dE�y,f�,-#�}[����(^������@��p���&0�;�s���wq�^��vN\{�H�
�_cA`�p��X��B���ϭ��^�	uɲ��TdS�́矘���ڗ���
��}m��m<9*3	���
�H2j$ă3p@e`(�>�NK����5�|)��pi13������ �OQ��4ղ �Ytfw�Qf�ڝ��sU�M2����$�A.1�b�ʫc����# F�5�� ��X�]B������ <����������@v��w����iK�0�@�����A�� )�J���<ї�6jDK���Pg?���1~!��W�:z��8a�5{x���<�0�`��~��k��g��<~�G�O�%�)+�������Ú{:�#�n'?�X�<��������r!%	/��`4���F�"<�6r��:�~��@x�un�k�8uO�Sn$\�^z7!�6��+���
�ʥ\d��6�^Ds�Z/����(�'���L`S�:E)?�`��8�'�Ā�>�1�gbݛ��6�V��2h>b�6�n�aC����7��H7U1�>��+VIU�0��Q��>U��y�s���}�*l������Q�[��߅P�ƋA�k(�z��*�����Z�3��̲5��Z(�T���]��~� �"��+����+u:ہ�%Ҹ黰�R��_'�=\҅���T0�����Lη#��]@�����d�(��1�G^��X�h�93X�7�;�����G�[|���`~���T�t������c�R*�~y��<���X\�¹3�Ώ��d1 ���)��T��Qd0=�� ��w�e	0�`�7�(]�&�5%[i�tTQ��ދNK�h���7��K���BkE�q�t���i���:AC������;�YW!V�^��k�yy���F���M��~dO~�%,Bf��7\A��y<f�^� �K�x�Oe:>����?����^�B�
zum�i$�P%8$�r��$R���n����6_Lb+��I��B��>~.۱>O�q�@*tz��H���|M�5�_�N�6?c-v�D�(g�4F���Z�2���(Q^��L5��\�XK{�� ֋���x,* ӿG��~����dN�8/z��I�i��%�*�!7Cbo�޺�gd������͈�\^#G�ԩ��v!�h�A�G7F?�?�n��-�n}J�Wl��w�	N)L9Od��M�FIm��*fn�Ϋ�����
����"�+E�RJ��/�e��R�O�~�����D��{����!����o�i�Gi�)��c��Ǒ��`���	�Wx�̆�7����Y��~���	��b`�s}��~���=���bc�ł��vGn��Q<�>�]�����dp�a�=#�Ď|�Fi￻���2���H��x:�L}t���&���{��+�~��$ɬ�li��ϗ)DT��If5�4�hyAt��:��u�N.�s<�f��{I2x$8:�����o��#e��ĩ�;^o�G$N�Fj ��a���ٚ�oi�(W4�蝤2웙�Y��H��{c�3υ��a����0Im������
Р�d�v�ݝE®ˇ�ҩ�X:0��wÞBpPBɷ?;w�u�iT��7����i�^qE!��z�L���q%��@�'���9+X�� ۝�����E�>��v��x
���N�̗;_��E�M�d��;��m3I�ɔ؂V,q�C��~V��3�Ы����/W�ʤގ�+�-n6N���x�&��
MNP��6oܐ Y���v�f�KM����+�8��t��-1���Vt�o�ڹ)��;a�'7&z��Y�D�{�E%B��If��x�A��"��{��Pf���v�}��|����P.
ء�T%�v������7�N�Ic��k�@�����`io���-���u��KL�͂i:�9QD��k�c���ׯ���2��GxiBm�R��˕pc2�Q2�˥�s�*̜ȗU-��/n�^�w�6����U�.�)�W���p�嬨�e�m+��0
	N�l��]����`с7����B��ﲮtL���Յ+�|�5?�s܋΂뗟^�a@n=�-. l+|x��F?�$��ъ�a���!�>.�J�m� �����d<� j(��)g�D�Tzo�P�]�AO���up4�`�����,�O%���5KBn��8��9'vj�p6C�t�
�߀D.���d���$��{bI����Qˊ'��ҳ�(f��>�EB�Б
��*��bbd��>Z��-�1�!�X�nIv����S�ƙ��L>�9ͤ�`� �[��lt�0_5���.�&:���q`��&�|j�������ƹe[~����p��cf�-r����`Y�6�g!mh��C�O|��ls�?7�j��I�ЪOx*\\�*�,�؁�i����(iaفຬ�˹ ��Н��'�d5eݛB�!��]z��1'��S�9y=Wf�ߖ����x�^ː�Z���S/�� �݋��W�uŸ�F �Aہ��B�t;�Ae�s�-�Ax��[J�!�����0���>��T0��A��Q���e.^�-	�(У�{�~By5�1Il��L� �������X���\Np*�����{��؊�j�s�zV%�H���|D���4�cxn� �F� �3�}�lD���JY�Zq�Ĝ?�%��H��f�`G� ��꿟U�C�E�b�!��fUt�N�>D^�d��'��\~�#4���=�����6�Sp��.�&5�;�'kݸ>=��z6�Q�2'�u�Vhݴ�x�D��z;�%3���ZWHi�.����v�{�˫:��W2��f���]'������X!R�j�'2�0h�I��q��(wG��N:�<v��+T֤Y%���:����S1Լ<�|�Zm��K����@S2�v"T��*gt��w�ɼ�o�e-})bC
�n�ؿ�{o���R �2`<�d�E�<�B�ȝbP"�@*�D��y8+�!�FRrV��h���\}O��>^-X��$�:�{�W��P�a� ���fH:y�A�$?x�
��6��m 45������7�f�����#�a��|���(�8G�O���E�z������X�t'`Ή����Xp²�2�
:.�Is
�����?4kyk��������I�Ɍ�<�9�w�?m;ejD�Y�R��4���1�ꝛ~�(]�k� �S=*�m��Y��ro�M����$�G�Zl�fȜ�ю>�ǥ|"IP!��Ʀ5�Mt�\<)*m1EF��n��$Dn����&.*�e��<�����KUh'��Ǩ-$iH�ȃ�m��;�+����e��n;z�<܊
a7��&=��+�-��Y�}7�]C�\W@�^
W���4ԳO0p|!��C��|gL(:Y��
�b���=%�<���_�#+�4�YZW�/���2�Lb�܉��)H��H'Of�W.(���I�G�[nՊ6����|�����{���,������V��r��� v/k����n�a�3Ql��v��yNC�KJ}Y�\}��>��7��;�7������OT47���MR� ��ض-:�n9=�l嗾<�W)�G���{E�+���Q�oC"��ylX����eU`�[�e��k�ӕ���!64��	"�6q��!�3�F��c��)�y�K��%D8�Į*$m����,Z���a<����>�`���lh����8�nu�����.ték�ȉ�=3jf��7���0Y�ɺ%2_�x2JQj�&���c��#�/���,*�,�b^Dn;w=�����Y�$~4o�&����?y�9%��H�m�\����yRso�Ϸ}�;����&Vn+��!m�[������ʞ����݇��e��	@i;�8�6�����[7-�$M��pW1s��SX�W"�D����#�ؿI�>�Ⰻi~P��"O_OVy�X3���Z�7Dh�41���N@{x��p��� ���!�k��ӆ�aP��
��|n������݉��=!B�s^µ�F��n�=9��ez��:PF�P�=�Z��N�?�;f�'W0ZE���H��R�yP���Y#�P�
but�@lh������*##�4�?�o]+4g �����*cx�@]c_%��S^'�i���1��k�k(L]�%�j��Ml�RȬ��ZǲKt��vk^�賣P�Վ��]�e�6�T�y��1�>O"**�q�G��J���PY�c�͔�����AC����M��<��\��R0!{���4W��
��;d�8V�-	�T��nOq�d+{Đ=I����Yܕ�R5�MhK$���ʠH�`R��[�R�CYw�_�b� %"����ݾ]gd�^x��@π�Ld�a@��F��hD��Ñc��Gy@%�õ�@@�$��o�I<���",136m�~��=�<y�3�1���R��&�=Ѳ|�?�ea�}���)�1��_�t;8�rP�#^�w�zx� V`�w89���7� ��A�Ռ�Lԍ��� �m-n���q
z�:V˚A�\�2��O���[��=�kJ��g߹A�S�.�V�b�_�����Mr�D�������-)d����Xpe1e�@����Vj�h@���^k׬�(���?�c��	�z(c��+t4�,�h-����2�Ԝ�ȍ1����I�ۖ9%�w�n�������$�&6{�e�;���+K�C˃��vN���Q��n�
���6�G��n��3�I����w'GET���Ir�h���mj1�ƽL�]��wP�KH�r� n�x�̜gnuQ�N��6���!R�Hi�2��p�O�m��7�/�-"������n����=� CP���+�����ܻ�^�M\�Q4���B�E~��ͯ<	A#�%*+�`lD�C�/�6���s3�������6��2A���o�n��E�|�	��\�P
����p�`
V��H;� eJ�'x��&��ʍT�i�XiǄ�갊"�щL�y��d<\+�'��=��v�3�8�ek�&�L̀?�Ԥ���6�nG�8��Z���d\�Z3��@�t�_� >k��kz���Vs35��_H ��\�b���)��̘o"��wT�皽��Y!�`C�*��C"���:�.4�KȬ�{}�8 Tª�į�=�&��_@��D֠l''u ��L0|���Y|!�Zy���e-�����ط?�W)�v��r�5�<.D��@D�_(\�s�*�Zꉝ��tHV�SИ��s ,H�;"Øe);F>�ǔxt�Iع�սc��L`gr)��Ayj������i���L�(���z��@1m0={x�DM�ً�X-�8q}�ilf�K��} &��-k��v^X��UR��Plu�)yH��Rr��o.�QX��S��4����dڬ��Q:aw��)E���*���%|D�LQ���U���yb�W��ix�3m_爂��2�Uϊ?r��%�St.��IV�MO��i�Ly������El*����������Ay�Պ �a
�nJ�4��nb9�4�@��E�e\i#�I���f9&�x��:Y@-���M%2������+�x
f���:��Q�l��Aԇ;%������ī`��=*�&*܁cI�t����E��D~o���ѓ���V((%�1������I�c�A���Uʥ��?>��6=i*d:S�b]�
�u�7#�]׼G��.��TJ�|����]�w�)��k��ݛEh���^,'��X�2~Qp�7_�.�O���(h3,�V�B%7^�e܁%��<B��Wz�ƀx��~y�X~/�p̶����zWib+�;�$\0���֏*Qw��&���\u5���ˁ��� ^ pT�@z9�K*>�[��}�OjfZ�'�1.k�� Ԃ���� �=a��e �Z8)�b��	?Ȇ��T nN��:ߠ>��
�'W�@=9h��˩E㧧0>e�
#�)��3{̾�$��O �l�Q�L�a�|Ӊ�$����
����nńF��j�uyʐ2	\��8�i*�&��wE	��v��L���?�EC���+G��Y ��)���Qu=e?l���[/j\~��9w�VV��8�����ϰ��:�=��߻��F�}������z6��M��V=]�/ �}�I.s@�Oy�I�ߢ(�����<���I��2_!��{������Y��l8p���sXcU��w��p���q�����Ł�.��<@�s
/ޞ��d�?�+V�6�lӏ�e����� ��ݸd3�ڨ��h���#Kg{K�	Mym�%ա#./�!�$�ϰ�Œcsٟ����M���wSdQ"��5��!�./t�p_5̀ ��������k�i�%x�C��޺�l����M�|Y=
T.}]��3��6槿�bG�l�� K�ľr"�s2Χw�X{d��'��)|�R��%?��gt��C�&����I�h��B���
�m2Z^X�,�H`���8�aբa'P�Z���'/$��i.j��#oO`�t�*M �:�,�*o�FJ&!a�c�Zą���7��y����B1_�.|��W���?�,5'gl�baE�v�r/�X/��M���v�r�dN�ʺ�H���RHL�����ƚ�%�����S*���[�X�%R��et�����<s�Rq���CU��3��f�Hw{��#�`1�<G�$���r@�̲٦��o!3R���#�m:'�[��
SxhSi��W 5l�/`H>0?n��l�ӭDe9ct'B�q��t��Na�̩հ5����q�\���M�!�"L<-q�jq���ֶ\�Tb��Hp d�͕�W�QJ#�K]l�l����!���6��[<��)q��!�*KW�c\!�m����WƘM��r�ǯ]�8�8�,����@�{�쀦�r�kC�������G����"���~�Y6FV����C�,��x�g�DwSE���@&�nb� -��fi��~	�]~���+&��@v�]�0��[���˝K�	A�
�]�U!��t��*s�z�kk���*\�=@�fY����P�!��J�w/���].��K�]��$������:c�PY�ub���Ӭ�B9�>�R�ʿ�6$߷�?NW�,B�s����ٟ'v�
�`�����P;��|�<ҔY!5A@�<��Gv��׼\-��֫4i%���^��6��V��0��$5�ӌ�o݀^��-ڈL>Ad�6U���&�E�:;��q��$\��fף��Jj�6�̙�F�˒J��w�!�^(�,cr�d ���E��U��x�5c*8?��s�Ǧ&ߎ*Kf���GcX�Ѻ�����M#��H�T~����=��t�k�Y�MiD��m�п�=x����%ٸ�!.�+ox�o@�5Y�4
���)d�+��PT��*��[&�2�:[�F�,�s���,W�l��s�d)���.�HG\+{9:q��s�=0l�|��Z�U���r>�O�?"8q�z����N)�ΚCq # ��}��>�(@[�)�/�vtD�8�������1���oS�,�ho�ʧ�V�K�'A9H��l����2�� ��M��j��\���k �a���#���\�o��1:G�T=?��� 
��gz�e�< q���_��VQmZ)S�R���L�z�*���Iuj�^sZ\����/�a{o��iMV�}&�	x<�7�քc߳��;�ڥSZ։@��O��@�C`�}L&��2��4y�-����r�(G�N7LM�(>��g/^�U�{Lo�V���-�:C�h�x�:�^H񙣻m}�J���3�c����D\B��>�н���i
�c5I�H�	'���w笈mq#L{���%�h�Q^�k/�<�Pưu�)��o�<N�W�3;���2�_��%��]*�˃��U�U?P*}�,���%�k�R�����YF�� 
��J�+
q����Z�H�}�7l6_����8a���z��F��o]v�EA�O�w�4�"�a�ks-�� �tfܰj��Ƃ۱�z%*gA|����`���K��v�����}��Il�`���wA�_�xv��7@������|:��Z�?����@�,T#�k�����!���5�ǆ�b��	۱�+�q�zӍ}^ć���/�=be��t�]���8T&U��Kٷ`3���#w�L��g;��_M�ܑa�@�m�'��������[�S�zĊy�I�QL��sG���:�(�H*x_'r��7��Sl�:���ϑ�� 9}Y����ioY�nѪ�F��L[����@f~'��~Y��NNm�j�x2�E��������e9�,a͂B�u�v�ěҍ+"4���%���� ��sy(P���˭�-��U���T� ��s.��+���5F��&WK;��j !9�E�;l]��3��	��d9��-���Y�cF����#�bؿ�N� X�QQ���#�X����-���8i� ��G��?��:��c��J[i�=I�<�3%[�MǓ�#j^U�����!��Wg��~o�8����B!�F�V��0u�^-�nQ2���lc���9��PS��g�\=����V��F��!3"3�?��|��{��9#�r���d��'�6�j�H�&�2m�ғ%����+��1�QH��?�������J8n8|�� ��$���S��[]�mv�R�����p���nk�%�����	|�+�&�E�΋Bcƛ�(I���4�$�$� I��S4�"�(��o#�MU���z�'+u�ch>3�q������f��x�jܴǬ=b�	J�(��Ǝ����D׀s-��IT��C��^�ѩ�x��5������Ǖ!�O*��� o���*�w+D�:Ř�W���q����Z)��M(�۪{�[��N%Y��X"��[PN����R�"��=�n%�뾷X?�-�Tۈ�)���Zm����n}�-$�o��</�F�9����M�A0t#���$z���A� �BT�ʹ�-ʁ��<���a9Z�)	'���8qk�b�F��É�X~��66�[��O��e��&a�J�uRʸؾ5BFo~!U�]��med�D�N�������.S}Ф�8���=yTO�����lh���#/J�cXBP�d�xb���u����@����BJ��g���G~K߷�^<���;;�G���x�
��{e��~Mx���7i9��tRPg)[�&�峏T}�r��,Dvu���N�J�~�Y
�-.�R�uD7�1Ŵ���T'��w��f�v5������z���Ū$;��N���w�0��-׮�vJ_����'�^bL݆h�GU��Ƙ�']`Bo��j'=Z���s	5�ԒB�;	�X�4�yo�:�r��a8��Ȫn|�\=Bm�h�=�~�A0��΍l�LHG/�����xKt�Z�>t5�^|�(�R�!���I2V�e�O)��Z*��*�������]
u����LV�Bw~�	KӲ8?:�U3��W  Vk��1ȥ�� �����6�}OAv&l�N�RQ�Ps-���N�	�7��=N��a`E��<(�j���+-�}-�!���iX�Ȱ$�G��
��z��J�Zƪl�S u���s]qZ�]RgL�I�� >��wΪC�4��fp�\Ưyd��5�!�"?�	�yI���F!�^MR�6���+��p�I��iP+N���B�Qy3���S�f������M��;����[���_��p^#�p� �:oA�u��Is����ˌ���CL�E�<s7�6#fɿ�I����.'�2�a�O>oJ�/mw�hqVd��[��:UBaO�誺V}����L&�2O慪"�o���H��ɫ���=xr��2x5W%�lD�M*������{'�nJ�>S�ש"����Ie;�rP�l��2�YTu!nl���&Qřȭ|=r������%XZL+��?cU�P�d�2�x$���!J�E7�s?�����l�.���\d"?{�ZՀ[F��6�Z9�/�޼� ,�[.���,l�+����l����e���թѹ'f~�<���r�� g�&�|���*-5R��Q̋���K���v)V�\ԡ46_tQ�]��s��4�����!
��J�O�~�Ps\�xZ�ck|��h�1��n^	~�����4��%0��k��^"��ݥ�h/5�qݾ!���j��j6�
'\OHr��hKncF��j����倡v�xuY�1��*v䒢�����~;ƴȣ3�<�7��j��)�#�s��t�.�Vp'�S����+o�X';n�烲Ɔ8��w���޾
����	`��P2���5%3dꂙ19Hw������X�U���rf'E��C"7��9ʉ`��*�̠%ڮ���E"�P�ֱ}��7�,����8k���c4ُ�ٽ1xp*���D�2<B>�l���"��B��P�o�j٭c�-��P�M����}k=GI�8U�[��_G���k�[C��H^ym�]Z]��-�cqflG��`-�_�T����c������+̊�³ �c��
���#�����1��M�s~�Y��<�Iu�;�:vVmX=!?4�n�b�1�c§IY�'�kU�	|M5��}$�|	����Z5p��q7{���z-�����ހ�3�q�������v�ֲ��SF�6o�$��^�H��ax��G��.�Z����(S�c��D����ǔP��GV0Wd3<�AIo�`�n	�>���l�������w���lU.T]<q��)�<y��B�m�R���yJ���S�`4�i?|ң#��,�P� L+�áu����r�S�/55DګAWnv���A�[ �>D-�My��APs�����R,Z��OL�TJ);b4�چU���鎇�-9*��o�[�:l�wyKWI;$�ڟSE:"��L��=�YC� z����k��a��W��+�	~���4���IE.�h/W�/Jy� �s#��riW���������9k��x��3[*H��V��6R[T�~_wO:Ϥ^,�~�d�=���W���N��)P�/�L�ح�����lf7�������nT��!5u�탳�`Gr\1�O�C]�f�[oK�1��`�`�F��"\�\W�Ը"?�[+s���i7Q�-��1Ũ��m��E�|F�ɱf�=Ս�Jzse�}D��P�%d��Z��\ $T��S�-f���d>��ea�m&��؜'�C���4�kn3h5��;sVZ��ɇ⦽ 	�y���ق:t�y@����*=����V'�Yk�w�RF�>���}� ��Z�[3�����x��
MB���Rx��\�ͩo����EĕA�[���Du�;cG]�j����&(O&�7�s*��-y�-Z��0+�����MH:��h����~ 7Il���M��,�_r�\��{, �xx.Hc�A:��0���s/��,ܖiN1� Xl_��R��Dk��aF�A\@�9��Ocr�f��9�'���#$WlP 1%���Zb�W�X��*�e)��Oˢ#�,��w�9�2����'�Ï��u���6*L���I��	����,ZAT�Y'H\1y�Z���*��"0�P�W-K>��M�|����B��0�h��wɪ1��l�k^z@��-6E�%'?�q�o'���70����|�W��2����P���ˉ[Rk�H��̮la| �nL�B5�������'�6�G�`�u&5ta%����7	��t��yOy��En����k/l���.�<��V����b��t�*0
Q�ٻ^��[�֪���>Ɏɴ����ѳ�����Fi�yM�Z�w�dAp����C)KS� ��Qî_gG��������A�Di=m���>R�a��r޹�h��n(�u�򬢖��=W-�v�ƅz��sy�+��_��^�֜�	�+R�<T5d�;j�� ]�{p��5~R��eD�ܞ��sx=�c^%�n4��?�b�Uċ �F�E�fF/�G���$ڔ>U�=Y�Y̭*�.��ZAd��,�D��g��L�v",�@���c�}} �0I!Z|B���-�v��?��J�Q\Zؓ�D㞡u9�k�Z  &�	�l����՞�\��t���y]��oZ�ڹ��}a=d+-�5S����R|���L5�m<7;d��.oH�fK�����n#�kىj�e�R�\s�%�y�:L��ԥ�"8��@8J�7�R+��`�m+=�I����m�@���7��˥�B�tI��7�C9}S�R�j�h
�6^ ��uf8D�7��+�a}QI�:�<����I9N1p�	�{G����x�U�i�����Y���^!`�8D�/%Dt{j��F����~�);��)aik�Kw��ץ�&��[;��{B�A����=wg�@vﺑ���n�|X����ڻ,����a��F�,p�%��/A�ke<2��|�J��`6,K��k�z���P�|�6	���yB����.Owc�k��^��v�eU2�M�ܿ��Yz�&�n{=u���n��|J��N٤�iv�a������qr+��e��
���U�J8��X����j�G-���4�H3x�x݀��._O��acu.}}��ɿ�'��폑T0L5Y+E�{a�A�� $OƗ��-vԵ�(U���A˜u�e��F�[���~1V���E�t������u��C��$���*�c������n�����R�3�l%u�&DZ�z�%6 ���"DvҞ�+]�mb�:��-w����z�0��V� ���9��s�Ft4ʎE��l�p���"Ϋ�� ��c�ӷ�́���%��"'J�㐰�+�B��t@�q�G�#�zKZ�G~5�I�vQ%�v0�
�:r�y���c;*U?�`B��ɧ��<`�9��=�߃��O*�Hg���H�~]�8���Q��y+�HK��p>��%j:8	V��?�+Uo 2�Q:�fY*B�{_8�i|=���4hYԘ��E58:Dgxi�4p���P(Y?��ɲ���&�u@$�"�^�f��B�3�JGu��̰�ݱ@���d���_;��!�q��� �ޞߞ�Θ$���)Ys�����ʰ�ػ�~z<��Ą���kI��U�#�F�O��7�:�Y�9��d�bby��>��R�%�H!!��vG����P���2[�<�V~=�]e
�P�e`��qɀF%��A��|*?����# ·t�ߎ+�<��a����WF H�q\	��!z*ƣ}�Z6{
�
㣀�nb�_i������}�be*'�¦
.��[�n��.�8=* }���-�$����F�}G���+��̆� l�.�m��!��>�h�=�y�D�| ����zNDi�'vk�\�ZSӧ8�F?}����)���ѯ���~4Z��˃�~^W�Թ��L\��2�4	�ܝ�o�|�KNIO*7O�'�"t��R������]h��(���!���0�����I�&.z��"$�;����3Q؄/���骇W|,ݟY�?�UY |�>���:���K�cr=���V�׽$�C�"�ʈ]��D��|��Ǒ��N��b@ঈEԣ-��l�[�J�]휳W����;���9xq�y@љ�i�~�k�_7��.Y,�,����EM�L/��_W��8�6.RN��_�W+�1�� o��4���_h��#2�wV$��mc����i�x崝�t4�^�)�&�2���J�䲊���X>J}ġ���ܶ��"Q�|���U��)����G\�\�~<W�Bt�ZY����9��/��:*L�9��5ft���Ε7�۱L;���y�tT�e�1����;oORv��E�C��L�0"J��hH
�[|�|���`��4�[�,8�G�M�TѰ�F��_�_�:|��06��M�v��)�\�4�yr��9��<Y+*O{�΍-�u���X9�aTFJR�'k��G�l����+��ш!`�ZV�ׁ�E~��`F�<�h�6��(�ǎ(Q&�>�`�	曏=3 �H��W6���cϩ�NE��v���eu�6 ��`�����h�����[�c��\.�"��*l�afi��Y���̘hi	&�Ʋ�S?�~ �a��jh�=6d˭�W�����Y%#�!��4t��o�����p&E���R����zI��y���$� R#Bt�
	��[�`ϴjx?�
Y�KG�[�c��	��/'�e�T� )L)��"2&
g���w�Ip�5�H�YB����!�ً���av\ͺ�����(W�yH|H'�*]����1G~�� ��H�Hثr��Tj�I��vS�������lM�DIu%���oLt�^���s���F[F�=R���Q������A_U@|sp�O��H�v+�A����6�Շ�_�7���
�	F��W�	�I䓠=�,puA~*�Hw�|�!Y��X�S����۶tO�������"qtw��&���0R^�	b���l�LQ�Ix�l@eե�+�@���Ǒo�R�*�d�����	�qt�;�LB��(�����'�̢ ���(�!ލ��#$����"�2�y��1�#Hi�zS����b��#��J͕䵃 hܻ����E�e���PA��}D:Z��be�\�y��}�}�)�����;N����v�̙�������B}�h�? m��At����1�r>{*��$'���nD�&����L��}BIP�'P�ցCH�V����q"�E�f˖@p=�|8U�{~ץm�s:8�y�`!���g���F�j���Qh�sWm�,1f��q�m9��dH���q"�j@��0+a���蛣�A�� A˾W昐BL� �	[�ǹ��G�saW��bF��iv����  1�!NVZ���S��,���FW�/��?�J3�80��SmE�CC5��T��&jo��ۢE~N���6�R`����AT���	OKr���P����L��f�76���F��@�S>��/u�ғ��9�}�Wb2����� �y�MQ/�-`hp�	'���h9��AE���A��e0�<	�F���	�<E���?��jb+��ӿ�P�(�\�͟�1��l�}�͚^�u��j��(ϝݾ��da�l�G�(I˾��Wr����L����X�4 ��k9�V̫ͯ��m�ݜP4�K
�Ԍ��ﴉ�O��nl?#��\���%q��4F�����-^��G���?�������s�����M(��=�oб5����":������>�%�U�C�,�?��y�֬��.o+�S=,�7GAw2�M4��c5�h�xA�/�Me���_��8{��G`�{��eF�`t�l�>P�!\!,mP'�$�y��<���f�ec�7�P��������f�⟛2�#�vʉ=֟b�9c1sx�*~��V�=o���'/Oǀj���D�C:������������U��ݧd��W�"o�}Ї|R����e-\�� wCO�Z)zHm��sx�lے�q�� l�߂�%����@�ʓ]�W����K�XwNU���F>F�q�ͺ�Zc�$��ݍ��In8d�G�ו�W	���Bc|xY���<��[#Uy��o���q��^S�G��6��q�+γ�h�e�u�<���5��J�Gs�b?�3�Q�LE�9�V�l�]��<�
	�į�אUT���h��-��	"��a�!ӯh��{Q�M��n�6~#�����z�&�s���b�3%8���m���;Q|>���ҕ|�l�IH���zK�K]TR5�H:6��)TZ,I?t���W�Z���|���k�ԛN-���+���r49'�"�{pbW:z�<��e�[�	m}�e_�2����Sݱ�~��I��^'�偈oK٨~�礅����'��!���4?}�z�Z��׼g�i���JԌ����i)���{�����J�Q��3 �5�ࡰ�dT��-�M�-PKp�E��n���H>˄7*	��AţF.zP�>d�C��ka�>|�JK�D* %�"����z����|�W������#;_c�uү��D*�t��yB�P-�S������С�6ǹ�pw��}�v�&���
����j,�n���T|���ү���܃���">N��LQq�a�qN�0}�cMg�,���W����t��`7G���ɣ�RLy:�'B`�꭫�S\�г~T��ir�a�<��*]���<��;X����m���k�2_**��B#��� ���#�mb?��m�PFWz��|�g��Y��m�W�fJ^�d��� ��@��Α�z�O�/q��a`?����s�u����Sթz���9B�.���P���V�]v�#E&��	�I���l�)�jS䟀X�%%c���"X3��X^0����?a��<��d�0��Ђ���e�(�91v]�H��
N�F�����0|fxZ��W�\^��K0�mf��k����8��6C��j�ehLi��#��v�x�o��:��*���ԆͲt��ۙ�h��t_�d��t�{Krr�Y
s)>�U�W���{F�DHK�rx�A�/ ���L�[ 6�e}�+j�\j��+��}S�Y��ݨO��~'?*�?4�k�^�ʁU���G�p�ο�, ���h�+[|@d�?�Gi���w���lte� ��pq��P�'��z
�T\4p�>�b'�IoK��Ȣ����|���(e$v�ua�PB�����vC/��cJ���Beܚ�x�e�n��'D�(b)�2��-�Ѫ\�}}�m-{]���C��ƽ|�El֚[�o:c�d4KכI{ȥ9���}e0ס�8�6严��8R�+~�$w�Vf���\Z[��us=|�92&���O2��?�qd�1%%)޴?����m�"~���4�gV%M��S뺶��	�6�o_��fLF��@J~"?KQ6�B\[c�K5�żMl:��g_�a_`�O���5�@��R��bR���a�1��-�w�O�����fT�$'kI�X+�6c���]�f<|7��ab�X�[V��9pWfʡ�C��\�����uw/E�תp�E<Z���A���n��|(��8�����R���X��ж��lj$D=�
?��uK��ϯ45μ�w�4���AluFU?�e*��Y+�<�l�=���Ǚ!�w Z�<5���eț�5Ǥ(�����	 [> ���s�ԥ4��k�KQY�i-?��ݬP��\ޭ��]G��N�Ʊ3�Ԗ+J02�q�lq�N�Y~#L�FǶs�d*B��$;�g�0�~
!)n9l���[�c��O�شy�[p�Fr�E䚶U�@`O���2�u�7(IR+�ݳ?s�����ӏ��%����0R���0�T�냵�q�AY����C �@��PQi~]� s�o?ۈˠ���PҜ�.V��D�3��>��b%>)rm����oo�(+��O{�E�6�qK�$Z��.Y+b�T8�o�'�ҿ�d��4N�\���/�l�T���= |���ɵx:�}�j���.�����G08���ȴ�OuH@����k�u�.I ��5��}-�,��v� M:n�h@M����DSb�jj�'0������A)�R�M?��Ӿ޸�`�t�1K����Uc�(�����@���>�׵�õ�I9�٘��i�e���	"�����56ƺ��c�rd�V0I���t���ƠB��S�����g�@:C�����B�(��&��r����b����
�a44��H��I���е(*���D�>C��[�Ɵ����{AeP�WV�̻�	���T�_��D]�H�S(���`����J��=d��\
���s����\�� S�ZZ�9t�H��)^�usCI�N`sD5i�W����wK�:���r�1!��LG��Z��+oBv���zX����i@U��k�3��|�{����x�{��HI��l�� 9J�"���K�zT�p�򞻗Q�H�z��ꦲ׸$�^;F�LN�p���j�񯒭+�f����tt�:K�W�[di䘨�Xf��V�^t��?X{z�U]����7w靮�(1-,��H�UQ��mǨ��R��lE�< �]�iw���#i�_�jݎ@�Ng���q˿�5��Ȟ��"��!�f��x�P|��?�ꨠоs���.RV1޵��Aڡr+M��}( �Ԇ�=���D�֜t�Q����=s\9��n��!=#.
����8���"�o~���"�`��
��Otǁ�r$�]�U��!Y�>,��^�7���B������Ť$�LS�*�!�hI�ԧG8z"8U"�A��Q���C:�d ��Z�Z\r?[/Lz��a!Q<�� !x �ARUxh
����B���DV��6���7��������1?�v!zW=w��^��Nȏr��?�"pTRR$i��T!���tP�f�K�gj��x����s����xʹ�q7����%�?��ZS���Q�{/ĉ<.m�k�X�މoYB�bk��@,�	*��|��o���a��Db��j��Ѿ�26Z�7�RRp�z-r��"Jbh������D�C'��P�zS'��u��^ݣ�C�:�{(�Ls0o\��0JC���ٝ���������ة��=�~�c�p���)��y�2i�nрͽ%��!{9vI���Wa��M������ ���2��t�]�r&��`�� �h���9ܜ! z_��Q��Đk65���tc���97t7�e�x��*$��0�ٸ���-�;����ܖ�m�w�v�`d!C]��je�.�o�וz�gD��:8�`%�i�<[�4o7B.���b����"��&�{b��B}��72͑�{�>��iT4���_�^D��^����K��}�8��2�~Kg�|��ő�>m�pZg|��(\->{��N�#����<���5�5&��F�PF����� �	;ϙxtx�)4�o�í��?�&��՘ca���i�������\&J<4��ٖ9Z�h	L%9�P��LlkW�,׼��n���뿝�B:��K��`��i��а}��m��F��_o�f#���Ѹs��%����x�xo�жq�CG�R�C>ޔ��{ S�<�@�F��AQ$�&�!�g"���Ј�ϳ'�wR���*��(��V�Yq��he:m9��/Wȷ�t�n���h�`�����7��+�]�F��63hc�Ϧ��Cs��~/@�~-.(	7�������8��
C(w�0��:��-��M���T�c)�YV��o �3�1���P����$����.?b	O�H3���1m���
�	v�ڍ��x��-^�d�"���pVJ�6��=S�.������O��l]_��R�����:�F�"F���e*�|���NS�8-����~i�;�I^��Ӑn���+p"�)������K���&c�1ܚb1��i(�� ��oo��֭���������)����E0��9�l����[��x6/��ǆ�ki��5��8�����,25mj�C��W��LYec���'�JHqNw�E�d.r�i��6�`�!8�@��Dw�6w��Y����I�Z%.����K�h�q/b�Y�Ŋ�:݄OG~Y�T��WWQ��(����#��X8���HZ������ð������	[�<��s-�& �j�h��c���!�?m{*��q[e�zhd�t�j���%T�9 2 g,�MQ$n�R��O��)K��-���m^B�$�|���-#�~ӝv�Fc$��lX��D;O���d r�3�d��س����>�tͲ����L\�6�*�<��t������y�vPkX��$1�;���O�X�����#�7r�4~(1���`�k��]���]��9��b`��Z#��\a��`w��3vݙ~�m���A}�0��{��s���zk�I].�l+��r.�1*5���B�G�9")�⶙��o�0��}4v!���B�EC��H���~�my��q#n�X��pB�j8\��{HRR��m5�6�G" �,��C�|�����3� x�b@uU�Q,'�X�y�#V��=������ཱིxDn�@��>h���i�zܴ_+c$�~K�(��^��nJ��/�M��nh�	,\��E��N/�\>�!Eu�,���!�A�2��~�'����ո�gp)� ��VZ}��g����a4�vV�u����T��%��K��M�+��ar�1��b�#=�2���Ar�	T;eO��eTG}���2�sd'��-��h�o�V)b�y������JVZ�@�r���	LˣEs��|�/ǲxa �]�$#�ƭk�Y�7@6d���A���/�#<�l�`�fp���ޒi��h�G?���'&��q���Ka�eH��*�������*�����V'�Wjkd��Z���z�oW_�݄�.�M���r�)FlXz��9��K�&c��]q_�If,.�7�J&������&O4�������z�"��r����F�{�c��f�f�j@�E�:�x��:c'��%ʊ@�{�>A-�:{m��YO�d�{3�_$���SHt\ؒ�9A�����<W��&.�,��ٔh�O�xj,��ZCQ��e�cxI2>'AfhW�C��*2��x��%]�X�a(j��߯�ͬp"@i��������G�fm\l��j�`��
�<�*f�A\��	l�:��LabB'�l��`4��o=�<Q���s�+��S&��/�8���mZ/w�㯺,��r{��\1�b�	�V��p��|��.�0�q�+� ��W��ݥOJ�X"���:ss�J���b�)P�͓:	�0���/#�J� oM�,G'3��Z�!\v�D�eV�/-C�=��٧�~�94���U����y����䴊�25�<�ȱw��k�w���������������� w�y�~��mH3u��a�Q�?S�(;��[q�H}vr���,I8Fpi:�X�+lpM��7}ȤLҼO\������c�kwa��/��i۴��T
u�����<�U�C�Y$� 8�2��!޻	�F�r�QH{����0�]i~�5II� ����Cj����]�p�z���ޙVן�qǴ8_K�O6�<����N�
͖�n�s��A�$$��;E~z:H'0�V�A/C�E� x �b�����v�)|���h�?{�|@uS��02Y�X�S��A���i�^r�Z�푣o�H='�?�Z�լY�㒡%h�&Y��^�t,��/�$/37�[h5��y�`��e����KW7���nG1=��pUa4>�+�e�,��4�T�߭
-�'�G�w�10����n�I��T�U��Cکd����ۓ1�¿��W��|��~[!�`Z�5��n��Yب4ԄF�_��}Z5��5M����V�$�+� ���ǳj����W��v]>���l���֢ɖaM:�R#�}i���_a>���J'�����+�5����mP� ��L�?)�T�B��T�`�၂��5��e��=�ַ����z��:m�σ�%����A\GI��8[�]�z<��g{�R�`��*o�
��/��&�<~�	�Nv/vU������M�. ^��D'@v�B�y�ƥ�3���XNF��:����Ot��.�/��;nms�8�mѺ�*dSTvŚbtI���?�
?] �=�Q����v�_�[u0��1d��l�c�d��R�HZ�����::��fx�d-�x����$aG���~]GŔ�UJ�V<I�˭���kXÆ��D)�� ��C�S�/ϑ����NɛyF��?RK���0��9�(9x���xɶ�[�ItA�%��E��X����T0U�b����&Im����B
y��JZ^1Bϫl���:~��)۪��O��A��2*f���2B%$��5���iL���zw_�Q�9ݨ˩\����:*X�5�1
�袵�����v}aF�JV�]��\��V��b�����Ң9�ð{۶*���`���p�8MY���z�s	.�_IR7������E�ӓ�R���A�EʰU��?@��,�l2�x�q�ztr��I`$���끅8�m�޽螙	<5�R�i�`f
���[�Zbr�~����^#����L����|$��k������mV1e]_�9$��tfe#�c�C�E܆D�v{��~,2{�ԍ��O�GK�5��L��V�4��*9����M=�����q��wv�	������Ȟ�� ��������1�w��tٽ[�b��EK��Ȋ�
�Uiν�ҹO>/n�з��N��HgDz�sscP,u'���v����*k���k6~V20P��v�W!�M>�?������Mza}$Ќ��g(j<��<9���q���5��Z���}��n�XͿ��,��M��nDM�3&^�Nã�����6��p�����̪j�l��Q���f���9�0�p�.굺５"���/��Iy��/J5�r�bA}pEZ�\�z8�\Az��[����Z	���[� �Lz�
I`��Q!� ��7n]��Z�����i��f���Uqv�I�g�ya�T�':$�	��x�.E���Et��v���}�]�r� �AIa�tmA)�yAxJ��F�!c�R�2ϩ6��A(�{SJ��l�"�[k|�Mڷ;����XO��i���c@]���n��Gy�#��t����;y���Ì�I�i�>�h��u˜L��#[b�Z�"봕ɣݴJN�a�Pw4d/1 �WK��N�RfK]Vg�	�Ā�/mn8`�V�Ø�=���y�mv��Ҙ7�EwS�R�A�O��u�� 6���Y����PzK���d��c�^/�N����h2=��w�b��:��4ǟ��qO9�Q�<|L���G�x}��H������7����l��R*,�t���R<V�pǤY4,!a��l�Hl�S�x;�,��Җ�A�
$ȕ�mqn��B�;��t����P��#u��	wEw��^laa��%�7��pmpś�2҅�7\���d��"�B!��bM^��ӫ���o�B�d 9
@�iz4|�E�y�4>X�RJ������H����@�}g\!���D���u�YKܘҵ�&Z�0��.y ��{����om�;�OE:� MՍg��H���a���QֵD��2����
M le�9i���iT��?Y>a���O�Nb\&3�p�[�V���_�]w��p�xw��la*U"�G��@�eSr8�nﶶl��Ÿ�+~%a�I���;�N��#ci��g�����Im�y	���[)�9����V��̚&<E5׃�c�p느?h��u��`������Q���Z
���t�|Bf8q>a��Z`�x�S� �v�	�㥒x��tⷍ�'WS�~ۨ��щH�J�ϔ�)R���(3P��RF�W٨��vE^	+@V5� ���X'���,56@2iC�t�{U��p�ӵ�4ߚ���T��K>DB>� ���&4.zv�A��ʍ{��͋����n(u{�nIm]�N��<K��1M��F���Պ����ϔ>�7a��T)n�l�$�x��;��E��?�Ja�Č�P�j�?���裀�B��k�!��I�}�G�4x����̑�צ���0x;Y;b`˪������T��9S�o�/�1���aFfp�;T��nt�7C�U�F�a���C�$�-�"9Dm�N���VV����dV�R��k���Q���*
�
��NUw,4��6S�D��O� �?����~���=�e��F�k�f�����b1OOź����Z�C�Y ��G���_N>{�=�>]�ˠ�|��N��l�.�rmru2�0�+6�->�^E�H:�2uH�7����0�^��"�.�&c{�,�k��܀b~$+t�I@q<�e#��To��]4[5�^��s�B�x��o��q�1�S�.��+���I���(�)�
�p9�"�S4A�Z�\$5����%�5a̾}Ӟ���ɔH�B��+��?�I�}��
�^|���F��Y� I�^��$KC�@h���Sǖ�s�S��7��'}�z$)ba2'��C�@X��7�[�OY�zM�oάT������Q?̡�n��}��X.%;��ƥ[�/�z0#i�'b����� Y���Ē�v&��EPy��;>L�X�S��ܳ���)��}��)�K��@:̨J�-����dl��� ��fY��S�{̑/vv�g	�ۖ{�^�Iu�����O϶N�r��U���ȠL����J�$�b]���t�y<���4���5L.DL�S�4)7`�Zzbބ4���}���W�R���Π��ڼ6ת[��9(��؏�Rc4a|v�ǔf��S�������$>���a�U�"�2�3���+�Ko��������G���5�@�x���_�b#i/�&)�((���@@���i�qbw�f�:#��WN���VÑhf�I�ɍ���s�έ��B@��@,)D���޺�~����B%fd����U��켣U%�������:!�����i\��e��ky��ĝ���#�\���������M�*�d� �r�����T��m��s.D�Õbx"����{���xp��(���B������<G�+(f�����zS�}�?�k�&��V�Ζ����sg��<����I������{r����~�����K;� �u_h�	~�>٬���g��p��ҍ�d�C��!��J1�B:�K�B��U���(��*n`0GP��I?dG�9�s����<�:F�r�ct��]=�\t��p qf���2��%L�T�˧�7#��*��0,8 �\�, );1Ϧ���cK���SU�8K���o�PX�!ߧ|�T��_��et��nwW�A��Ԯ��/������dXX2��DEO�a<�1�ט��;�俌��T-KaE�@ؕb̨�?�Up�����jĴ�������\_<����cC&�Ξ�s�S���ű���ܕO�����nevd�L������a��4�.�]`7�N�ĭbA�6hGϻF�\�[�x��E<s���j���/��}�*�<2�K�[h��D�wɜ"Qbh��3���J˘ ���X2�'�m�j��G��^��C��A��=�h�����[�K+����I ��M��M�O���>�:�
�ʿ�=Є^��&!r����:rZ�58�116��ܝ�z�w�t>,a�\�s��rƄ'b�t�\1�mP}�|�a(��}'���ۘY �`��]%���=2�S&��6��r7���" ;Np,��_r��ym�:
he�|m��R4L*����?Щ�(��+	|�N��=N��0���F)�:R{�u�� 9V��G.�/��l=K 4��m�~1?ٍuU�l�5����+��XtY8P�Z���h�s��	��kc9�0��fj�2�Զ�1��ga��~��J���.�+5%R�d^N�^��頡�0S�`Ǚ�M_/E�e�Î�m�W�y@'MlOΠIwg� J�ꈹIN�1�\���]X'Ogs�ȧ��>"�_���։՟���ؠ����>�1Z�Q�L�����?彜�2��5F�B��J�>=�Э�'�㉢#�vs�abǘ=��t!�|����M���I��=�G�� ̓Z��5�
���׵k��^�~qm���^�v�(`�k��.4Z`nU���;��'���_����¤y^�O�VCwe
?}^҈��Ku�?����T�֒�fɴ�i>�cs�xp��ߐVTe���ߩFu�4[)��[�bu��n��`�B�<p�0��J^�6�Ir��	�YΥ0��D�C�/Q�ݭeYBo7}з��Q����܀a�wVb������㨷�zv��jg4��#t��EVj�`!�}l87��l�b"��I��AC�
g�B��G��PS(3l�,�C��,�
,�O��i�]���޶����
%�X��gVRPa@\����o�͔Js�Ź:�=��)���Y&������i��*���a��mM۽ıU6#E�?>c C��}��=aٴ4]( ��<w�/�H��wչ���*!��(�!�%$� <>]-������Tȶ>��-��*hmT|q�
��%.5B�Nx��S���HbP�e�s���	 ���[�>kC��4�/����Y����?��K�Nf^\j�i[mE����,�:G4z�ռ[���1׃C���׏.bq��C�-�^���VdԼ�W�Ϻ�X~ڌt�1h������;+H��0��A6l�}�m�ؾ�G��;e�4���6���.X�$ %�id<T�3�J�]�k��#�B�;�nͻgi�f��ɧ8?�p������澳3���˨�@�y
��)�&]�����+��Nd���K0�>�3l�+'�'���<��x�BhL)��Ou����p,�=�cw�9���߹��T��!�2�Z������D���@����m�Y��5c֚�'���V3�$�n���>�P���{�L(���ЌǏ�\Ͳ�k"���q*���L��ciR:����.0�ޘ 3� 9BpOos��t�<��̥�wR�D�7k�)���0�|�+\������'�%���k��~��0G�{�Z���SB���l��� kph��7��$;d}��b�&�9^D#��+C�K<��H:tch�j~;gx)�o	L�a��
B�ң��^��`�ԑ��l��ZH�L���0��VU�Zz���5�ka`�kmg����@�B^fQX��ݶ~��`��,(�&���=����ko���=��	F�#Z5�}�LB¼;;��\���Dv�qDz�Q���ֶ�]h����!�j�e�ֆ���1��?��K����~�r��/�������1�D����-�"�fH�)��E���� ��3ӡ��ᄞ+A�G�`]c�xG��f���%�Ӝ�>�N��EA�=�4�� ���ˇ�O/��f�IX�;Z�#īZ�_6�v�asJq�Y��%�����d8�|�q��f�._b��/�B�aK�O¹�:��~�C�6Knr��\ت�l��,<'�;:4f����^���Ӣ4O�M��hwE�3��o�N�g���^��P��c�pfq�ch:�E�j�#7��-g��dB���lmF'v��pƞ4��	߁T$O���0��;dǷ'��>J������!����D�񩌀B�Iy]���E6�㇉��=	[w|9µ2<.Usiu8�ۺ�!|�M�dv��?���7�-����f��k9��W\�qL;�K��i��ڨNaZ;u�2if��ɔ/h��X'�^�������Z��dt��"�8�߮$=�'�J��7ж��]1��pxqK�����Q��0Kn?�s��|2$/#B-U:�M�sr�_��2�Œ1���z���E|ʇ�P:A���,\1�B��ɲϰ� IZK\�.�߱^^ ��4�9H(����qP��D�e}�T�2o���,1P{�	�yc�����(��<�2u���XhvvbB�c�5.�x�l��9cg���'�!��?����e.	 S2�,���oh���7���4c&��z��N������=X�	���\�])���! �]��e�Kf��@!�"�!uMF�Zo�پ͸&t-n��G�3Ӿ��t���7�������VR��ڒh��Ƿn{�%NI�l5��2�?3�	�}̧a�'$v�k�Y
v����k;]�%o+��������}+����Y��q|���#���w�%�Đtq��ֿ���*�,�۩�x]����$�	=T�O)���뼑?֭zȋ��6A��^��Ƣ��f�IQ�qL�-�x41��<�e��\�;CLNr:ױ�d}N���*���	w��V�jԻv��Xk;�����b�ͭ�%D@�&���3���Ő;�`�зߺ�E���ɥ��j�n�}#.�
�vD�Ռ��bDN;"�V�Kbm�9.���"����fsk�HI0v�����s�crDN4�1mLY���1���v����UShf�c�>Y�<֘�m�0�f����C����sʦ�l ��Tv��a�ku7��� �9�[k?@_"M\՞:����Je��!8��yld$.�� �O���h��1���t�ۺ6:G����k}����	 �tT�nyK���_�!�U��1dC���V����C��I�uD��n�U!�c)'7˾��0�A�H�ѴY��4/�v#�I�䛓��.¬TE�r�m���O�#�w�V�w.���a��X��c�%s���#+�JAD�㵫Ԓ5�c�-�TI+MW�	��>���PM\u�w>e��̂Ǒ�$��B�*�&���f 1)�� i�C|>ijL�"L|�W�Ϊix�0���Eƣ51k�-�8fz.�y�E?t�k�1��£A��8h�m�T����^	t�a��sG��C������NR����"f�$~"߿S�3�'쎺��6���C�\�W����_�"�l5
��|��"���Q���urM�ޢԢ*43U�%��q�9������vv��Q�H߈ޮ[̡�{��|�A���&����%�,���0צ m�	g�c���ac���	���̝V�Bgh�|.�h8Jla�f��-I��d�� ��m>��M9w�$ҁ��eɺR���Ꮸ�$�g���:8�h'p3����֯u�;c�E�X��R��1H�â�I.9sS8��m����xSD5���ı>�k�y"Ţ"U-c��f)�U���]>
�yq�Il�_r��A�\yJ�~/eR!SL	�sW6ϒ�R}����k�B���	��I+j��9A^>��=�t���/?�,�#��~�@U�F-���>�~m0��Ƭ�m�y�?L�B��,5���IX^W��a�$3h5Yo,`)O���|��)sK��\�����r�/��~u\	���[�29���w�]OlG�jt]��_�M�W ]�1�^CyEƅY?�;�C¶L�<(�T&����xqkY��1/�s�ƒ|4�{XN��D(*��ꀰo�x��N	��v�2�!��N������!���
vAG]��p"��	�F8r'�D�� ��`�/o7W��&9j��c�Ҭ"vh��(!�D�b�Y|�[K����Vɶ�z�Z�G���4�[@�L5���9>�ߝ.��?&v���V�Bx��| Z?��Q��Q�¦�~8���kGP�x�ߊK��=>�?��̉>}8��#�!�b���+����	�Q �	��T�xrpYЁ]Tu�	���JJi��u�˛N�v��sq�6����~X[PA� Xj�1�L�hx�w���i_|�#ag������`��q�w#D8�j}��\W�$&I�7�Pv��d��
D�تv�|��d����E��*�O8��)���qP�O���Ihp�hI��Dxl@�1���f���EP+,���ʕ��{�w�I�5$�b�Ί1�ߤ�Hg\ٚ��]���p��;��M�>Yk��:��Unʈ^9�-���(0 x�7�0���D�*���d�X�1;t��;���f��((>bL��>�t��>�9)�cT�?|���yȂ��?t �;��quq�l]�Fm3B���g4@�� �U�dCG�9Y�/���b�ťi����@Zv�X���R���q�I�0�����G��ꅇf�v�<��\�M�t�'�S�o�U�?w/�.���>s�~7��Ǽ�<�HuG����%�Bv��<�Ԣ���٣;��@J��
���K�{�#/���|񴧷y���B]��XS���D���7�,��&�MM��Q� � �-i��EM�ew�ݡ�2� �:˘�Ơ�@s~W��K|�U�J�(����F��gQ�FD41��&d� Y I����N�jN���.I��at'85"(��O�t���[���+�@���Dj��G�Z�(�t��U�#",szoR0yYs�9��jF8��!gi�ɒ�K.���< E��5t���x�����d�)Tfa�S�7��4���	���6h����-8�UR#��ߚYҖܭ?�*X#H�s?�� ̃G�qsowg�#��/���-j1ع'� �W�~����*��nɆ�u~�|�L����<�A��n�a8$��k|2
۲�5��s`��wF�
��B��a�N� Ǳ��N�1��5̞r��d��f�¡���<�AO?��W� �amZp�.��R�x]��pӇꪵ��N��.Jӆdvڈg� [���X1��A�$��a7�Z΀e�[�{�+�Q��v���R�����]I��k9~2�_6�Fb"E�a4 �YW���4�H$w ��,u\�E��]ǡ��M��`(���߼�OX�1g�M�#��2בֿ���h.{�(�\_J��u%̞���*�� �^v�9|�A�YVY�]�`�D�9��Ń�����=,�^���Y.Q�	����~k�ɱ�R��4� x�����yl�]�Z�}a(��ۛ��:����,u��`'�!�q���Қ�5�O�u*Yhĵa@/�	e�݂�>v:?���f�  �6�u�SP�M����^(�����5��Xk^%zOH�K��������}ԃ�_�5��VJY64 �/��S�>"��-�ف�l��P�=�C���ԑ"Y�Ӓb�n����'L��"��ɋ0u1�5X�q	a�Ա�]y��#��H��I����츲�F�yE���*�v;��L����@���@at��!�^ѿ|��P�=ͽ7L�AZ .�+>aX=�&+JR���^��6���X�w)'���|�JH���f1D�k��kZ�����ô�)�����Jw�QV�r=%Gc�u��������l��q?yP���τ]�%HXY ��L��6%�x��lup�r�>�y�@+���T�ӯ:d�%R�K�Q�e�Z��`Zg����N(�5��\���%��u���:hn�z���b�G�d��S�F��%�ۊ�E4�ͭ��r��
Lo�*%��ݶ0THѕ�]��#�Ӷ�6��}`zd�)-��U�Az�mܪ���Z�FM����Z����C���)b�]��+��^��:��N׏ٱ�^w�4��7�`ap�QC�=�
W�Î�o���pZ66��2�v�(�a������N�_�~��˖�@����V�JK��z��k�J�W
��	�����
xt3n}��!׮)u?����g񶯹�{r�y"s�]���A�vQ�M�v�XK.���bڕ�3�"�?A@?Ni��/�1�7U��ֲ}�ս���薠�;k=��/�IQ4��h٭�����R?M65���l������	5�������a�_s�� ����*w��=g/N�5�b[���o�u�>��%o����*ւ��I�;�PS�+�>�f�smr9>���Q��D�ˤ��.�wÀ�0�UpٹW?�����r&��z�	��pU��j,B?�;�7D�9�o��LN$����1����+	�k�{�ҙ�d�Y��{-Q�v�ES�/�7)]�ÎQ�V�iWW�X��aQ���SH��v�,��Rz]Wã7Rf��Q��Ԅ��E�&��~(���Gw��o?4;�e�"�J����"���X�&������CIC������*Ak����\R�>EШ�6g�eX[ã��E��c-9ҵ�(I���<��?
׻@d�ä�@ۅ�$�׍��vڀ�j+��O42��i}�sw��sy���o0#M�G=����b�"�8�a�3����%����S�XOڳ�sN.^���V�`ִ{�2+Ȩ���0sq�y�2_�ޖ'G޾u�� KU	�T����
BԾ��;���9�
w�ػe�'��%���ۤ��j�~�.A���?�#� ���s���[j���j�)����^������%��ִ�̅�m-ۑw�"��_-��u��w��t�s��C�nʔ��Le��j/؀'A�6�0����sY�H�AR�{ެ���sVq�| )�zF.�>:KC����J�c|�A�~�fVl����-��1_��AA�f����xټ国�c�K8���Fa�Ԓ
�䗾(��sg�Җ�s+K<�O98y�;�Ŧ����٠��e\9���q�J����6�A�P	�ꥥ�m9�E12F���^K�!Q{��/]{�~vlu�E�x�B�$���.x'����s({�*�\��*s�E��
�U�� _J����f,��^�ra��+3���C���Z`F�c�elӺ�c�tӯ�F�OG���wH��N����<ߢ�����ٱ�Ń2G�@�����G3��?�sié���8����Z��K FO	*:�����B�?��½�t\"�����_<�IWw�DZt�ՊԔU�t���#�����/Q:�J���� s��k1��F�QI8�,BTm�=�R6���h�۵���9?Ǡ]���U��[��?)�h�O�v��@�EQ�v�}���\P��O��v;*�H�빈a��Q��4���E+a��7�M/�?C�SM�'lL�ܰ���"�w��i��4_-�J��t�ll�L}�v�U�nw�Y<[�z�=n��P�PXx�15���C�����>D� ��[#6W��<��C#j��n_D���i!L�%��d@	]�;֍�+���Y ��#Nu�|F������=��%���᱐�b����V�C��y�V�y�{���/vLM��:�3��?{[D���?p?���z7�8���ݰ��:��Lh�?V���u���5qH�,�i��[^`1eo�g��Vx�R,��˷ U8ڡag�@�LC��G�2��e��f(��X*�V�ـ��n�[(��,��'D~*�Gȷ��v�#6o7B_�g��F�qh���T �D�%	���~M�l�1����Мg��7][����?���B��{s����{�!ε�B�YE'�M���LC�KV��dQS�ɿ�
�
CcB��փ��'�K�󖰤�6���6�봠���"]߬s"h��T������q�L���W�����gv!��g[ajhΌtR`��r��0�69J(K(h�>�L����:"����1����Y"��@��7����j���X"9���6	3���6��Ǫ�����0]�W8�͒��J��e���5iib�r��xh�Z׵�i����ܮV��ً����D4ŧH�>?Li7�MV�����3�b���͘rٜ�+�+�S��� tKi��}<-�ĤQ��	�U���΍�F8�n[8?��!(�&� F�}��v뷿�!�������J�2 v��"�re�F/���s��jk)s�
R0e�ٵIl��kq��֐��dvk���p��%,�Ta�m�h���[?B�x.D���ł����O�"迊 ��JSL�e3vuC����@;�����f�0[B��<	�<�x��DQ㹻��"Oty�l0K�[���1Ĥ��^��E�D�IH�|�&���z��U��ݦ5>݀k5X7����4�i�N��3���f���?�� �K+���U2�)U�K@먔�3�cP�hhe�|	��\ĄA��ʊ�LXH���׾�v8q(Z���x<k���h���Ы ���>.�=��B��ȽVp^��5�:.��6|���bͅbݭ��	���QMt��(��U{]�d�VX~�1\�wr���Ԩ[�י�k���էƠ��m߅���Z.w���+��Ql�[�3T��ԧW����0�h����E�FkGy��,�>4t����b^a�d��ɚ�4,�~���T���F�M�zxX�$2��TM�����ɜ�ˏ#={������/E�8R<kb�O����w�����\������w�G�wC�}� Y.��$54a��`���b�x%y�D���Z1qL��0��U���qx��?$a����R�;�ݞ���C��OG+Do�ﰩ�o���}��5&A���8i�d�3�Y���F:�7��� k9��o0a��W�|�IunO+��D����N�F�I������������d)����-�{Sf����С�"�Rګ^q�]��z���hFq��	zxT�N˸I6��M��w�e#p.��F(��4y��J-)�)0��|8D��:���|�� R�ԓd5	���O���X��:�*���{�5�R���L]�8�wF{��!��@��y��A:�v]�t��t��iS�
83;Ga��i:��!C+~U� 1��#��+?��+�k��dn@��t����@��(a���C{���x�R?�Y�j�`5�����U��!����	,;���R:��4�pa�~	�h��f�M����E�J�%�[��{`�kֵ ��h�ֺO5��EKvu�����j��/�m�Ȍ���=\�/�-��l���z#�8��^�F���b�J[c�c=)ʌ� Bɏ)8�k*���[�T���s��G�"�$c�^z�����Y�]��t�9�1ܱͬ_V9[�­�q�t�=F���8;��H�8К�a"*ť�1L�&�� �j<�R��g�-�i;�+�"#cW�Od����]�"��s��y9��� ��|u^I�ӛ�<Fx�ˮ�m�U���$�+�wګj5��t�ez�&��xS�������g��C�%�
 �]bQ�j�4�8�q>@iIU��ƫ	��V��u����Q��Ѧ��o��7�q��N&��(M��ڐ��M(N����<��"EMO:���/3�]��LGX�L��ږ���i(ݱ�f�x��iz[��B��X�U;G�r1�.�o�,H�v��z/DB:R<X�$���*L6�����˾��q(y������>��N���������ac 0��"g���;�2��'�9|H�IQY��å�=����{��6%�3ث櫖X�Ф�.�J.�O��Y�e@N��X�[9�$���)����E��Kʢ���­��ͨP�:�MO�[����M�a��,/��bG�'8�/�s4��P\/m��B����t�����s�@'�S�\�Iҷ�B�_�c�^�V���KY��A�Vԏ�qB��kK����ҙ�V^�+��ݏ���=�ɢ1?iiG���_ˎA8(�d�[�"���U�DM1P�Ax]ܯz#��[4�ȧ����q%�,j���'1縗���
Q_����$��G��-}�����ZJ�6�-{肸��T����Re�%
C~�i9�p���1��Μ[��%��%郓fmՂd*t왗���5K�����'��а�(&-�}<FT[-����"_�UQ#�!f���{�|�PYl=ҏ]��PX��b��&����iJ)�j�~# q;���4�j��J�n�̪�@T+{����6�!���Y�F6i~y��D�����̌�ѣ4�6���0�z+�bM��|�Dp��|��v�Lj��D`�K ͍�Z��8?��GZ��&��2H�2��ɮտ!!չ���l-=���u�,֯��F4�U���T�"�|Pp����t�Uض�@aA�;���5�<��պ��@N.F�jF*n*�d]�6v,�kL��!�P���|7kÙ��9Do%;j})!11����@W��k���(#��[��vIm�!��*?e%['9�~��v(?V���"d����D�FѺԌ�v��n�
z���@�*F���댁�\��"U�i�}��^�A�/ �.�z��L�@v�N�xɝ��O��R(�֑�>*��H�+���S�8��l	V�Bt��Z 8�U���]�n���O.�A��5�@m�X�;9ֽ`H�\)OE�&e1$S��N���#��u놮�b��z����~���X)[<+���g%���9 ��"�ы�ŗv3I���L95��P[�ܕ��a�6�NM�=�����գ�	�[2HBe�:� �nx�}������έ���� ���l�rߏSSF���Q<�B�'7�Y�a���^6[�n�`;=B�x<Y���e�8��X,0�.|�*�YY�kC+�̷�좨ޗ��\���y���-Yg�=b�/NB�3�A��Lq��C�)���
���Y^KG��B%W6�x���!�$���Ѧ������~ѱi��9�(8�:�9�x�&v�]
�h8p������?��y�����	��%z��G�a�Ư��LMgvC{�&:�����OQ�h���g�徑����	я.��œ/Fu����
���kɣ��P��;I�]���؃p����ZJ
,ڻ��E!9����x�#�q�[PN=E��q��[�Ye0�zZ�T��p�mV�u��%t!��r������G������Ì�����q�|��i�i}#�i��8�&�!A�	pW�y��^_���`C+�Y�JN#2���{�'!������Im��h���2��Q�ۘn/�YG���
�S����A�p�; (!?�;�R2R��$pQZ"u!lds=Zu[����q��񩾛��Ϙb�H�k��u\�:��jj����ۢ5�^r
h�h~n�2x=c3��&���b�ت{��������_)4|���4����Z5���nh���f�B.�U���}����i-,m�+$�r�	7�y���n�~�� IzH�%����=�z�j�@��ۙ{M@w�i�<W���j�ٵT7��9]@��$��P������)	����M��������X��9��8�h@���J\���
��xKt�`F�d�c�$ ��1� �0��V[�'�5�Jx  ��a�l�IaC�0=���-�IX���B�7F��):�;�Cb���ug�+�ruBp��,fO��J��5�#���P%��[{�.Ľɠ��T/=��D��_#/y��@A�~�1��q�/Cc��[p)%֛M �i빣)-Kx�{�g�b!3��##��*"�Sr�	��nM!*��:�@�笅"�s+��.�?�����{��@�Ok�v�7n�t���Ɖ5Q:��~/�0bb"%*/�H�<��D5�Y�!2���Y�xt&b�G,�eX�$D�.HVכ��|�]� =x����{�Z
���b��̭s�n+�1�e�W�2�n�:�g��T�����8I(��߭Ɋϩ�+3#E2� �$j9�̋}eZ���6T�a�5M�3�I��<�e�=vW �nO+X0�M�mP��;Ζ}��#�ǐa��L3�r� EsY��,��u�g�Ln6��kl�޷@:�w�]�����H+#bG%�G�+b�3�#�zO��*^��Qڂ�������z���o@h=��@�P�o���DJc�B���5��u�%�j+y��!:t��~��&q
�Ut�+z��CTz(�@�Y*��u����Lc^I��f��u<\l����\�����{AK�a����	
�V��� 9� NOy ��Of�g� �=>��,��K��_?H[���c��*~���e_ҼFf!!�H��e"��`�B5��^ѰŪI�ԉg̼�<\56:�b���Js�-?ir��-+J�6�Q����
��֨��9�JV�)
Չ �i+#G�����i|������ �Ee�rE���	t<3�)ѵTӿue�;H�<g>2�?��6�%���K��0�B�/�"<�ht_�ԏu�����A�	q#�]ŀ�q�w�^c�+r���j#����"�	�u�?j�����X�8@w
q��IA����(�k�G���[k�sOڀ,�&�'��a��O�)ļ%���գ0�dI��m��0����@p'c���N��ĄI��1�Ï�V������!i)�r��7�c)��o�</s6�d&Nѯ�(# �<�IݦL�,���"��V��Bva���~�~�D�%F�H�}F�ƽ�M/g��v�r^�����)%a�ˋO��BVl�G{��1#�]��Qs;� �@�X��(MF�����.)I��9*АhB��Z+��2>/x	��6��c5"�_Ҹ=�J��x�U�!���WW�0�2e�ܩT�x���/�%����x/���B�������Fa�� cI�N��3�p�����E�EVX:k<�Ӓ&������"e^����mX��8u8�(�zHi���4�
����(��C��/��r�9�?m2Y��V�-�|\��B�C�SOK"�i
�R�>�
qЌ���i-w�&SU�&e�U[�:K��m�zV�IV���v��X�0w�V�+];��9;�H�c��Ա�u���W3�KP�{��21A����qu�I�ꮦIK[�Of�ޚD�)1�5�=�XCQvn��O���%��,�,$�Et��T�:l��>���{�-9GY�╪�8��)�I�3���b��T3(.��2�C{&L�LI��13���5����@�g�P�f,�#��}�Y��k�? ��qM��������H�eڰC�֙y`(�רh��ރv�
�9�3->�KFO]9�\/E��:��>��E̽~ �$5�����1����cnI�#�v��F�6��Y��a�)s$`�pud����oM����N�J�òc�u�/�C���C�y��ry���X�D����M�������>�g{\�0^��,X��#��*�or�r61#cI��H���I"%7���Ę��	��1ܧ�z�W�(�0�k����:]��O��%��^�2�����v�^I�y*S��EY����c��;ߡl�bjL��c��|� ��s�:���1�Q�o�}H�j��4$> 8�n�<�c��3TΒs���������B�S/�P��+�*τ�������;�w��?�ك�)���z�tW��	�[�FX�;�I��b	�#E��̇ͧ�֢�Ϫ�lW��\�|3�x9��[��-������n+�|:R�m��RΦ8�%��L��0O�LW�Mk�@s����-Vl�Ϗ�|LQ������q��(�D�H��������Ũ��3�4���'��:�u�L�1�/��T6�B}�O{N_���E��nJ<��,��l�{2^z�	��NiG�9���ac�wd�9�X��s���C�tX��\�B�D���{1!��c =�kv��
�V�s�}�[\��f���n}���������� �{BıY��9c����B�jR�ٴ�Mn��	�"���0��{���XېܙV��D�~C�#�AC�*#c[�i�MK$��?h�[���}���[���e�8�h	^I�;�#�8� �+T�Hփx�<�&GLq7�Ph�a�?;lf����S����$Ft��j'6s"� '�w�6x?D���1LBd�֚�h��zwe��B:����#��.蔋�H8�!;bz�S��4zy�����c�u�[>��#
���Cs<�1��3n?`*g�K�j��)E�N�.L=C�[}:®��.�Z�.]��*��꣍�HFkV������5��W��D宦DQ��[�	ZBݬ䗲�ǽ���ު@<ܯ\�!=�f�{�:q��MRF/ ���'ް�nt�r����D�n9Ex�!�kw�e��H8��v��U��t�~��m�p�Q	cf)�KGo"P�9��d)�yr+�(�UdbAТ�E|�w�XY͹���؍�|U�sb=M����F]"������DNon�g ��w
.��3e!�^����H,q����X�I����?�t��0���ݕzv�a~k�ʩ�|��([�($T������\��|�ܙ���}��e�V�V�������3+��gb�E ��}��1�-�f�T�8�g�zf;�����{�!�vo���"���z�{Y�ђb�
��=+Z�Q9=�yR%�G��V�Po�н�0��nh}qr���Hf&)H]� �a��	˥X���1{c��ҝ�=Ε�>�Y�A��S)�w7�M��
���H0��f�w���FbN��H]t��Qӂ�s�y_���9�(1E���7�\��8��ה~w�-�%��Oď���K+-*/���g�{Y�㠆'=��Sib�-8 �~t��I妷7rK�[�޵J$����a]�Zi|����dS�|��ҟ4��{\u�a��6 W�`B�yf2�˞EU�F��	�Kvq)<��{�������*0�M���éG��$�#	��<A���t�0�C��#�J�o�n//��Z	���hA �l��J�� rr�ol?{��U�B��U?��kff�T<4�F���Ր�oU���wSc�za�RxbϾ��@J�5��8�]���.O����%KH��m�-��e��N~z>�i� h��1x�]:��HN�Y���b�$��'>SͶ�f�ԟ:uk�w�<����(]M��8�?����f-[|���
��P�z�pxgT�wϏ�ko�&G��~E�e��Ђ�R]��>l�դ.m<���EX��;g�� t�����3_�L�v������צ��'*'~��ѡ�˟Ľg@�'�g֒�O�-���#jQ2���@����=ľ�C���{��V��5�=�O��V��?)��`���1��6���wU"��<���ghBH|��~_�{/]
���*�$��/�?J���u������Ks�	y���e_X��,y=������*���;Vk�(É�o�oW���b�6��%��{� BH���^�Bm�K:8�B����7�M���>)����5e��n��N��&�z�(z
������̿9u����+^΢��/֐ϣ2���
Ӑ7/=V�9N�t���R�f`>2H"�w��	���̨.ዣ%�>4cv�����4�q���&o�F��W��ء���	�:��٬݂���zK��ؘ���Jw;kqƛ�e2d���4�c�z��*[��!v�mTk��j �0���Я7Q�y��ײ[֒�Β�ƣ�\Y�豈�4,�Jc��1��C�����C|ŧ\Bɿ���Y��y��qV&�u���ݫ:�%m�����c��ѣ��T�4t�SPR�; L|�,2��]��s_/�ϓ5���<* 3��d,`j�6������z.��o�C����=� �ޑI��nGA(����] ��h��W^,����6?~���yB�ē���Q�EЌ��h��AY}��⿚�vV��_uh2�FfX4��3%������ !y�ۢ�Q"��p=7��8bu+��O `ޑI����?T6�)�L�.�	���g�xC�����ܒ���E$��X�~$A�+��;h^���J�6��ŷ�.��P�c2e"��жL�.슝7���q���`��!�^���aj����􎵲���4��l�M�ue���8�Ɏnw�
c�=���}|*�a�3jR����²�8�͑]`�/ b�����F��vԻ�|;�!�bT���D�m#����s�qwq�|��f
��f�U�Wtq�9f�{����MnI����?36\�i|rО��P6�����e�&�,�!�ڌ8�M���I "1L%�*ʂxþ�Hh~[�t�Y�Q�?��w��bְ%Aw������z�׫5h�Fd�`R!#5��,I��r���g�jW��pG�K
�J�o���"��Y�����j_�%� �(J1f��_c�?l��S����o#��7�?��Np3�<w��b�T��Wi�^����A�T�U���3�V������J���$���gi<@{u�>Sa�)mȤgL�)�K�Qӻ/��xc	l�=�b�\V:^l�@�e�g��x͞��M�u��i���
{�����^�M�a�ٙ�2�i+��+��p�a)Q�4g�f�O{�9���L�;���^��m� �r2y�h��׺�!dqD������kX.�J�'�g�xr1��V�pZ�k���A�L���$>	>
��֣��֠��>�@�u��hu�J�EJ~��(P�ˆ�@C@]�\/*d����ĎɠYs��OggE�tU�*Zv�%)�p��[�Z��&�p�^���H��G� �@j���Ջ^���,XLgN�X�*�����XP$�c�z�[<:�i��xW�u�&ݜ�P�s4�֬Wъ���ʶw?7�M��%޼�^)yA�����V�H;�đ�U�5�Q�Ʊ�A�=j�Hs��k��п�?ܝ��2V�V:j�텵��kz����I�(�#I��2Ӏ8�B�蕈��nN2�ˡ�1bu�����vwB�n�3��Ib�U��|�&O�����⢅#����N{�uf�M�G�9iJ�|�D>���g�2�	�9\v���T'Y�E`:��7b�O�i������������� ���6����ZV��!e0��c�{�֥��|�ϭ����]&ݹa�%���7�����1h�%H�oCH0*�����]�  �'>gzg�Ű���D�X?�u(�^$�LA+���D�G�A����3�e���8�Q�Ҙ/�e`���ovK�����mZu������Y� Qp���Ek&~p}�89�!�S&�뵡�!���i4�,iIL4�+�N(����-�"��N�������\:D����Q.�f�����vt�;l�k��؂�F�Pq���syӽ& w��v�����FQھյ�\����9�0r_;T]m�M{��{�9�@�p-IW�(Z�gYČ�J�t�F����غi�RT��.�䄻�/Q�_0�ݯ�������p��[w_�`v��B���g�ے$z�������`���bN��J��D0Kr�+�/���%���y���wk�>K��h7�l��R�p�mc��L�Ghmk��^�GLmþ�F.�U��1�rc�)֯'�r��2*��`A$q����m�@�:an~@}�xvb'[Y}���Hw�&:�S5�ʑtIU^�"pڔ�&��� �����HN�#�AUKe����s�/��% ��ɷ�a�v��4�Z�� ��[{�Q����7��<ƣ�[�w,���H�1}��ml�a��;�ѻ�������ʃ����.<cɠ#�o����#�q}>a`�4/� �;1�Ú��Nܽjt�E�&|S[w��H��1�����޴�������"q�Il���F�}����p�ǚ�hF��]n߿�{�v܆<��͛w�Q� Zc
Xg�蝧����:�v12�9�B[�)��ql!٘�Cd��ы�Q��[�JM�C��^��=����WS�@�볫�6�4#���P"EK/<M��;���ܩ�E�)�8]mE��c)�nUF#F\c>��Ꮄ�R�M��q���Rw����є�Ɖ��q��N�}�h�p�����!�t���NN��̘z����19�RB����(�M��6��e�; ��W:@��J�$�Be��=�2�	zJ/$H��|�}l�~Y������c�2�>�)���-"o�<�9��u��z;䖄�[�2�^�䅍����$�,�r�|q3�&E��@K 0��T|��T�,ab���ݫ��!��>'�
�ؼ�k�~FU�(paUOϦ��L-&�n��ؘ��W'r�~D
�a�!�^��༡p���1�"KI��ZO�u�F3��f��i	n?�E��(�g����G�2�c�o��ZN~��1`:���D��z��{�)7ݟ���4��?I����;�{O�����hm�� v^g�$[�$|g�����P���e��G�VS���K�`Z':̐�*�H�[_h:w/�?�ޔ�4ΜkOh���s��v �����m]�+O�^1$�*�{M:h���'����Z�)�n��Ai6I���[��D08|�($�����$?������%�:!�q�=8��\?v/�v�gL�E(�ٜ��b���	PW��21�Y���15����A+y���
�t��"�h!�rq�B����Z��~j� ;���"������nu1(���]!4�[W Oc��!h`���+Z@���5��Z`��梚�/=��O���-?'x�\�t�"��zM�)������g�1������
���	��~^�P.�/�^H ��clM�W�|瘏���g!u���ئ��.)� �Ȑ����h�}2O�؞K����0*cK�NH�{(���0S�����9ui<3��*���k�lp�z^K?61��*��4�\��cH�V���5}]����F��4����TL1���SQ�b��@��旳�^t�Mv�Q}��(~�Π�I1
 ������Yc�G��{��^�ҟ�Z��t�]<��kJ'8�9������yb����?*��S�s+D�����]���<g�B�������;o]Q�h�z=-cs� �q�5��m0٧˪�M0$;����X{�2��M�}����|�4�Z���}S�)P��#�B���	`iWN�̜�Mߜ��9��-EP��, �'i6���MM��@�|l\�n���I�!|�kO�c��g����������x,O�urY�����68�Q�}���jY�8]*���q��C�G��a�E�����ųm�+�����4��Y��m�����.�5�B�O�~O����������ޓ�9�&��ke`3�^1��㠣����:(9e9��$ӗ�2�g��٤T���Ο���e�r�ƺr���/'��'��0�DC�|W�\\-ہ���=U��]
�:������	@�)��87٫(��a&Euϑe�lho��w�pktk̶|�6ζ�F'M���Lpl� &�%_�����a���d��n��,���Ĳ?l��Ƒ���JR��n3>�u��5����0f��[�*�5A,'0�:���@�w�,<�1YuR�1�
���|��i6g�ܧM��|�٢�D��������=u|�B=��s^�d�;��������qޏ� �����rjB��/8d����g����g��̼�VƩW��&��`���dY8�҄�J|j�e��VfM�P�}sk��|
47w�I7w�Q��9W���9Y=kD�δuhAN���� m2�u���}vj���R��l��7�&6�y�A:>*$���U[��F�/��l�X��s&�~�	�k<�^��ͥ��p�~T���6�#�_I�y��۝�.���\7?s8��$���/ce��3_<`~�I荝18)�G�����@�W��ӳ�l1O��`���"	_�BIkA�Az�凸�ԓ�ɏg/�k�xP5�1Y���@w��k�ip��(\�:�_�^ Zq4'oΉ�K�o��x�Z�ò��
���)*�VzFi7��y&[S�@�5HK{�F���6�1՛���bӉ�a*�4tv�!]�� ��/�z�{���v�6�^0Ԋ އy[��v�;�V�i΃`\��<���W߹҆��!3Њak;��<��/�'蒰8��&�U���מ}=��`�<���&��3��~��ezX�Z��v}�$FY�J�2�2O�Mab9����(=��<Lj�:Ku���J(�����6XH��Aq�SR�_��<W�hDM�����?d�V�l9@+Д{�K($��hߞ�$L ��ŏ{o�Ɯ�cR�����+��Sz�%+�}�p*�è!&4��g�Z�_��L0�e%����'���B�%餹��$�S���x�ا�p4ka���4��Դ4�IQ�Oյ\S����釪�'tp�|�x�2l΋,i�'�b���%U�J�$T��~��lkyfw0�p��+���kD8av��<$	�{�>�B�]I�P�)0d�gU����L9[�F��V��qN/�aP!!�J�&ͦ `^��sҐퟋ�Z�M'�m�T��̼��`��k���i�,!�P�IB��h��-j�
���Kh+8��1�Fk$	�<ؕfp�c�ؤ�6����G�i�Él�x�ܿ���y��e5;I@�ˉ�=��b�n��W���I���}�J��y��Ot�qG>�b�A6@-�5��5��a=��>'f<-{-И }�8i�b��%u{^��z1��Ցn�?�������+fbr��,���w�&�m%��S��<���r5�>��`�ueIQD����B����K���1�uE�؏ԉ����
[W᠃8@���'5P�H�������,���=C���SA�usN���KW��j�^9G�q���j�G�Dm�:����OH�-+�c
͚Qʁ�@%���@�S'��mĺ8\'��e��3b�7�p+4���ی�\K�5h�?����Y���[fɽ�2^��IB��Q�>��*[�_�� ����],���@Dx�%�Ԍ���:�����Z���$�'7�FqZt��â��ɬ[y�*��ao�XҀ�+!��iRa�,�[����߻l�\�k�s8D�({�A�O,������{�w�:�lg��xe�x1�a�����njY,������t<�	���U['ki�(6����fٙ��Y	7%NC���nS�қZ%�����9���=N�S�i�@3@9u�98��")pӵ:��W�Y��N\�7�����:�`G��\
����,��2	�W�XO���.|�E9���j�[��fuU`E�Mn�4�v����N����R�.r{��P�(92��Z�ٕ%�:	�A�i�ZP.^
����#��Jj��#�Pk�Ζ0h����,�g�;ū�������i��}�6�%oɄ�N.s��S1��?f�{���5���5�"nvb{ʕ~����t�0��)���K����;��*��Iư������q���c��tz{7ψ���r�j�[�.�u-��%pd}�,,	\�o���4�fS'�G�5�	��=Bu"�E��5>���6��eRb��v�̫�>G�>l9B��%|�ǋ��Z�*�6��H�&!�s�|u�$3F�4�Ҏ@��z,�:��N���H�2�ss<�jh\^+Ә&��$�p
�� �D�|�{oD�*���T�������G��Mk+-DE���֓��'�� �f�E��͛*�ZI��+�.)�~�>RZU	��P�Bψ���̞�]��r�Hε׋�[������F	�=q�ś�e�h�o���ґ9��8�X� \@
���|������:J��N�Vb��e轻�0p�s�<���Y	@��G��S9	L��X�Ɲb�~�Q���}T����f�=�Ou����C�б`v�֜��;�vgC���)%��^�@�\�+~��HHx�������<����`Z	��>#��h"|�q&�Jj0T�\�n��mnfD3��<�s��#� u���y�5K��>�P�u+�-5gu+c�&�E_�EEΟTW2�H��K|9�-��`,3g�U@N�4��dH^�ci�7 �':���S�b[�ј�5��ih�g⣐H�a
���E�Y�(O/ܻ���A��J�4�O�Ÿ�.��3�� {�@,�������[�Xܵ��F���1�`�	��S��Y!~�'�F/$��x���U��,�L��B�'�����{�[��6�GEd�p�?p{DV"SD|�Oe� ����
��L�Ea��²����
����v�y�����U�aE�§��������|��:a]� ���NWd l�"������~q[w�wba\��=4�����6+�������k}r\b�_�_��Z�����:��ir��{��1�Y}����/2�Fx}�^�@-�~��5K�R�;���i�xc�߲�˪a��Tm'��#�L\^�Yf�_#TB��Okx��K3�7	�`��;��F�h�F�-���vYta]Ez--JIK��߫�ۗW�ՠ�'Y}�_$-���!,��t��o�?nj9�*�}]Yb��)7$�7>�J�I
���D�g�,R�h�O��䡭�h��j;�{
�����
��}�� ���莓����No#�,�� K��^����~M�OF#�;&CD��ёʍ����F����?��0��M�!�Jp�w��r�g)dn�$��ޘ�)���l�������9�_�&(�FI�܂&w]��ڟ�c�"�9�����XAgDa!�3q�W��cPU��ݴNh���x��X��G�/RoR���oK�*��4(Z�C�e6fz���/�����-�q�xV�E�7�Eb�m�����ߜ�3�<J'S�t��
���])S��x��|q�r ��f�{h\wO��x 0�:����t�E�.��mt4�n��C�2�&!�ƃ�Ƽw$�. .'��5*]LџE��ĹVɮ����Ja
�ƌڱ�I;�-��x�m�X�%���8����egSr���ߋ���R�u�CR�x(>�6:3�e����B$�b<���n*y�K��hq�Qʒ��4Y	����	f���!��=�2�B��\��/��J���?�I�&a�0��1_�������	�泬U �N��9�7F�r�n^8��c���>�Kr�TR�^/�*�^���xS��3�I��%�J	 HGD�a��|yF�u��h7���jr�/vxi9�6�
f�l�,v�`tqW�<cѼu�N'u�=²J�J	�[�3���d���fd�'	��>$!�_ ���v�1��V���ވ����˴6��!� 8=���嚄 �ä|��s"vi��#҄�'=_�g��\]�v�k"9�V�d�����c�<E��V�����b��Sڂ��쿍g�<t�bD����?��B��}ad�VP�6"��V�%������z��D�T,%N��v�0�D���M^H$*:�z�:��̙����>���C�2�I�J��YRJ�a���2��҂(���'�4���� ���)�}�ڞӉ�/��_���k�����Z�+����s�������o�e:�
�����t��ZG4�x�T���	By[�뚍�1߷d��:��B�u���!��#+
cg�:�=�7�_93�ǜ#�Ǖ����	���;w)�5vr��e��62Q� �r	���RǓ\ڤ�]� �����?���eY&��I�!�!���,~@���:��u���z,E�)�Yl_�9�_�
�Ϭ�7���"�i4c��.�l��~?�u���a�K�u��yGEf4�l:�ވ�dj� U[u �}��>�6�:����ˌ��P�K���u�M���C�[Z#�p
�e�[ZZ/�}tU����������o��(�	%����r�B�^���=�3}������;d=t�,���^ncP��L���S��V49��o�ޕ��'b���+st1�d��
[���ye��
���o]�#{s�V<�d�:=y�k��y]����3��s�l���K�� x���<!b/Cr]&�y'��],Z�R=Ev%��S@�&b-�:oɏ�D
-���a'(%E.	'zx�H���u��^,��pg�Z���(���a��zNL7d8�їO��u��$�T�w`Z$f:(�&�(�HQ�<5 �:ΠC]q�Gh�b�ɺ_���6��[��ޣ��p@�M�aRT�?�M_6tD�$�m7d:�H�W��f�>��C��Į;�4�G� 
�Y�{O{%�J�0�&MPR4�f�蘪�L�<pJ�+P���`��~fUꈗ4�c�z�k��2lp��xǆ�u��1�N�3OMɠ*в�+E��
a{莮������Y�ES���(���`9�p(MSRJ���E�w��{0&�zGz�#���k�L����m�qG+ncsTfk1b��9�p?EO����je@�	�^.ՐO���T���I�N_�3li��?@��R^Ycj���/��P���ڄ�X��Q�}��6�����FZ*S������ Dy��X���F(t��VW����~�=�"j�&��L��//�ǫ�(���\V�|�G|s�Axh��;�hXχ� Բ��պS;1}N�م��h���-OI^Ҹ{u���d/ēXb�F|���p��o�r*��N0����T5�z�W)� ���@f�r��B�0l|���l�g�e�ē����8՟���
:I(�|9, X]��	?�ݺ�O?ՊЅ�[�S�۾��w�|�I���W(�߄��1��u�s/Z�6	*����(<�<ݲ���͈Pb+W�G ���=V=�Z� =�E��yø��Y��VP�}ȝ�g����L��q�ޤ��τ���q�ع��&�N��%�V���
~0�I���<,�����w�J���\�ڤC)E����(ӏ��.��=��#f�Y0`_<#rJ�
���R����:h��[�k������V���Urۖ��?�z�f�Emp�	%Y7&:<�ō�)�5`�����쟐�^�L�@�֘~)����3�a�L/�����5o�?�@��>�bx|���y5OЇ��m~lN�@$\�$HlPK��O��Ѡ���c�P��~�`��N��=G�&���@���S�Fҳτ������D]�m	��������Ϫn
��d�\x����C���P�z�\]��%��1X��ى��"��,=;�Y��C���'���4�wE�� �%���5ٍ]�.�M�l�`[U��������t������G���}�֒�2j2P�*��"���g�D9y������<������@��\q�Ɩ����	�?�����:��$�'�1zTSkxom&e�r�j���*�������J뼩�>l}���o��$ �X�<U	����V��>B��<PHV#ɦ����:��o����ǔ�Q��$��N�#�(e�E"���~��5G�\�r��ң�.��}��k�m*������@bm4��"m�M/�1�ZA,�L'8O�v�^#�&Q����n;N6��|��=q�B�<Lь�ɤ�`}����Jy�@��Ĝ��z�Jn9E�؛d�Ll�::%����)>1��.���Aڅ�\���"��x����	@�B�W�B�¸�s�����ҥQ��k(@ X�F�8'�xoqZ����"�s�&�O��i �����͒��a��9AE�ci�m ��u'�:Ry%j�~�i��nlľ�>G��u��MM��)^�\�ːdA�}i�Y����D-�Z!���i󥹶�^�SUpP�&�^��m-�!C4Ž�qը5�a �nv�%����g��6�n�f�]�a�o��ie�N�"�a{#+i2��@U܈�ĩ����Z@��ӻ.��3=�2k�.���T��qX�9ox�1�gY>f�fEL/�?�������-�����q�(H!\����T��B���K�,�ݑic���QV��kC=�$	M�Hھ��������ɽ��9pT~�N�0ЉZ����j�3�'}J����cנ d����Qjx6�L�nH���#�D*�i�%�0�H�`ޔ�hy�&�S�&�g�S��SR�%�_s�loa�Q�㤇(V.�������~>��"d���\�^������Pe�!Œ�l�Pv��R-�@?�MH�/k�H��7���W
��-W�1�8`e��U�S���3_����5	�W��g�I���M`M@HWf֟��w���Ů�`���Tt�<�u^Ƿ]x�b��+�Ȫ����<����'���ߤVEρ<�p5r���.|� �@�����ݛIf� *` .��������'���(��/��֬9_��rD**4'�����c_1f�i��$��zeL/Q�m�r;o<���v[��(�{�>�z@��s��gf�j�B\tb�i�>�BK� �G`K_��D?����c|�6�B�H�fi��Z��Ѣ]m��3�j�LO'{���'�3�����_+H���"<�.�>Hm4��w�
�B�Ŏ�C���{��p(��Z��%�T�*�I��1�;/��R�E����b!��g�ȱs�]�f�d������ �%��~�i��9�mփdu.�9������j��=��z�����mu���s��Բ\(��z��O!��}��^�7��K3��O��!@��L}B�8B��ON���fYu}�rX�%��Ӑ��T;NKH,D��/�Pad'���_��G��v�$*��Ē`h��$��r���FSL%���W�q5d�ن��NQb��9Q�Ss�T���*
s�I�ȕ�v�bR���%�Pqԛ~�M>4Y]i���^�Z%�� ��3�/�=!(ؑRPH�<��l�Z�w����L@RxZ�Ћ�{��_J3�z�!�Mage1�L�*X����]aȩtn�2e�I;��zu�z�fzH	�d6.*"-��=�T��"�^��U M$�������)�z����5%8+���@�a�m8�`&�۝�EV"O�7��o�o�#��KBbv�1Z�џ*}����1��V�����Q��jb��:/$q��߼�˨��g�o�(�T����o\ ��$Q�52O��db}��f6)%�Ľ���bG��"�6g�q�H�aH���ag 6��=�3��WY�\M��1.]������i���D,�S��9�%8��M�$s�
v@\l�~�z)��ǐ�H�c1�1�MQ{��F�~�7p=.�� �rn�P�a0�}�=�7�j4o9s���O�Ѓ$�.�D��4ly�Ovo��c����J���j��t���V�>�*�L��
���L9��7�O����z�$Wt��G���]7����B �/�ָS'�+����ԀT�!q�xH�`B�3��l��?C5�;�t*�~9;QmHR��l3-T�j2+9���N���TZֹ�����J��k^�i�r<TjHs�� H�.�i?�X��$�����Gf�� Z��F�o^��ՌT"�C�U�s��S��%�3'�<9����r��n�gx~v��t�r�:�ԁ�Y��ǔ��.9b��oJ�!ھ��e����c���s,��
����w@�l�ٱ^T�_�ɵ%���������g����	>
R���m����|�25��T�U��k�^�x#@9!��K�~ó@}���/�Gu����m�ָ��TtS����u&u��mљ	 � ��]�N�R��q`�Fӷ!�ڈ]x����Gc�ʷ��t�����B{�Y9�q�]ġ��!; [`QXGs�\a�X0�ڥ�]oJ��A�E�{|�+�Vd���{̶HU����HI��Eq�N���Mc�Ǆ:i9ԯ]��{�3�N�_��ˣ��X����#8<(�}���{7^�"I����"���^X�>��Ω�l�������Y���6�)�9���2�xM���I��rY*2Ha-D���Hg,N���5|Ɍſ`,�=�J�"�'LE�������VM`b�mؑܡ|H�ҵQ([��;nY	���t��({�d�^��A��yu�	�6����<y�[�;�c�=��|��6N�xs�}�=U�]JVI��=+���������Z0�����;d���h:����2j`l&�����<LX�tKc,�8��C���(@${�������u	H5���g�۹���d�ic$�pg_ӈ��As>��I�\��5�m�Qh���BE��q��959��|?�ۏSA����f��_��!�Y��9g&~:���;�kj�@J>/_�Hppd��?9w�b(v\F�ݯܗ�\% ��eo�$��%�!�Zl�ݨ�����O
D�V��5�����P.�;:.���E�V���okP��5�4or���
6��b��ݹkT[@���'4 �a�ը�򣨙������I;�߅Z��׹�1o�dЈ�Š �cx�����l<�aFw?�0��0��E����2{E���l�L2���[~Ab�QgW��u���lr����MIn@�s���"b���4��UU���ՙ��Ӈ��b��!���X!���9�l��W���$:!b��n�5�"m��@<DZ_��#К�g� BeG����~RJ$�:�̅?A�@�p7R���;ANL�PN�}M�2E��z7&m�|�\)�|a��� F��'�⚐��:gR��W3% ���4 !8�+8ռ�ʹ�aH���%t��	[������%^b�F�ᩍ���s�	�/����+��*�[�� �V����+:����^�g��Vc7g�A�gr.�Ih�T�jO��ojF!I}����;��@���\t9�c�d`����o=5_�p*^�U-q�z-��1�Mo��T��d&�kTƭM�D���y��B^��;T��,�����)O�fi��wh�U����:�_��n�A"��l��:i~���S��q�T�&l�'��ɸ�+�\#g�I�<�2�-:Fdr�������\�+U��a(�/��@ݩ,m�]����R-�γ�
Q#P��wp�t�b�Uq���vl_x�2D����$j��&w�W�h����p�{�;��oJR*{�eե���h0�#�N� 2�g��i�eov�y��@�ӟ�kQ�ς��`��}:�v�|��$J��x��r����/�p5���P>!��U�?��sn Ӕ֏�ܭ؉�[�KhD���|����tq��T��Q<d6����o�h��O�\��S*�Q��h�s}����s����(�{��â����yd&�U��Q����c�J�wk�p��vDt���X�C�;�Y,]�i�If!�0/�v�m3IA(}�a��A��A�)�̷���?�����g
Y�L�S�SBZ�7�胇���o�곅Ք�&^)��Ar#H� �%}� �UU�����jyQ�޺�E��E�b��+�?���5)&�~g�W}�"$E
��i3���&�y8!�=��C����/6Y�Կ�f<�����뼯CmD�>"������jK���e�G�2���1tx�'��L�z��t�1.�a]�����Q���x�&�iЈ��VU���O�?����+�0�P!�.�B
!���v>��H�è[n!@�<�G�h�N1��j�o��ᢧ�g������A-��h�|C��8�x��/��2�����*�LP��-�V�?.�d�~��ͪ�%�G�fȟLHC�(�Ց��PP|�:��,�޸���q��:�@X~����*ߠژ,������qx3��̸&�CQ�R-ن{�"�ᜓ��b�Y�>)��Ӎ��CVk��)�Y���-�E>�8�2*g��R�]ͫ���\�� ԇ��Q����DdvK;�Ja��5^_�W%��-Ϸ��Y�09�d� �7�J�CQ�{Nb��>�,��k�~�Ľ�ԡ���JI�g�;��l^����ZtM�����r�8p
�ϓp��[1*��#�{�Xya�m��U����-�m8y�r���9��_����:��GYl�+�Λ�\������|n�0_s7�J��$V{n��_n�2�'��Dez��#�F�t5�d1����qDdM^$[=J-���;?����~��Y��~���U���/�v���<a� ��e�`�Tl�Y��[�c��0��\��P�y��h��B$��sTu����=9�'.}�  ���n�ǵ�^&�^�(��P��P��)) ��n3g��ɕrj�-�ų�����Qrw�	������ܱ4��DAB<�oP�B`%� �}DK�%�@^�R0�n^��L0 3�ʰ���ׅ�:o3O�}�}|��ad����4�O�ȣ��p�UO�ѝ����:I���������~.��,��8W���y�-�����U�i��0r�[��Y}0�>N��`�.ƭ����)��Xa7w2��	U���П�(ȟ�|n;�����5
����r���g�R��$0
�܊]0�FNde����1�F������8���驼���F���m�&�Q�q�7J����Jj���M{t�ۆ2%�e�0)����o&>�#�L�������c`�f��9Χ��걻3<�P��Lύ�x�Ĭ�p'�E4���e,��ܖh9����W�lݜ���Զ�3��̅z��۪�YS���7gv�F81�q�]�oF�v)�y��ǌ�
�)9�#A�>>z�k��D����Ė�Z�n1��yEF=&�����lл��$m��Q� �M���+T,̄[��	�N���h�]fbLnW�h���aѽlY,�������!��H'�.1̎��V��6�:g�0i�ʈn4��w/��.�/�B{!X��̒��` �8pY9����d��8�W����b��i�M��Q�BʅI��8mzJ.|�i���W$5�b?[�«)*u�i�_��Q�!x��~^��"O�+��]��X�x6��^���h��J�V��͗M��u��#<�A� �7�۬�J�>q��z��	kxx�x�Jk������(���:�����6Ҷ�c�ӗ��J�D�����O��0ܣXtOi~-�*���������`p�n��\��D 5+�1t�7�������S)j����^͙ǯ&�m��W��P>ڻ��!N}�UNrS�L��F�Y ���zr��#h��i4D8�ݺf��w�E��Þ�� KN�0�
 ��#��6ӄ���-��}RAd�yìM���$~Na��֌���_g���L�5w�� h��āڪ�6�����n,���+~@`4d�.�|\%�q-R�O� /���s| �0N��1��{���Nf�v�O��gO�V:��d��,�%��m#�<mt�V������z��s l�m��[_MqC��t%�8Dey���Ď��\��#hMI�����F-� &?h���0�|<xA�J�d9K7�+>��t�ȥ�����3��Q�U�ë�����؁+����<���V��������`u�k�7��a-L9�o &�},�bĠ罌�T�����pئ�U$넖ʲ���.ޤ|�f��g-�k���E94����d��M�kb8�����>Y�uJ�nPF�K܏mt�Bz7s�\����N�?�9���E�A���e;F;:�=5��Id�iܟ�s�<'9m��h��l�����Pڄ��%��VQ�[㑀
���+í@V�X6��v�a�+�l���ڣB;��QT�ډ��wL"猡�<]U��eO�Ծ��bq�WFF�E5��E3룱 ���ʓ���?��X���M`�QHc�,{h�b��'/�̰�� `w����xۣKh����� ��ns
��n�n�b�0���D�j����*��W>��\;&~���n�O����Ȏ���v=9�,�o�l�AJ���ׅ?��%8mJ���&.�&���?g��sV����)ː�@SV���ӄGZ������{�$�����k��28�����j�����8.����cRM�/���3X�yd�~�ښ8�E51<��`bH��!�e���*��[�C�5eO�R<��������)ۼZY8=�M�Y�p�HʰdM���}S�`$��P�d��$�R��7r�s(���SN�O�om����o�9�F-#G8�0�tf}掏&˺?�-Y�!�9���2��Es�%���]6�&���.�]e��4��t��Sa,z1��$���( ��d�?�Zw�w6n�9HR~ea�u��{h؊v.M�h-a͉��R��i��YZ��A�W ����w�����_���1�n����`m�|��)Ջ���ڑ���P��Q�ٚ�I�� ktL�+�L�1��$q�`��� ��-�S��}Nbe�F^�Ԡ���#/�x��#�@�	#�#0�-��˱��^,�4Ox2��(�9i�V;�XJٸ�����- V���w씟(Dud�	�Z_l֝�o:0wa��xTu������V�� V�]��
n�Z�>���ZBU1?��e|�A�͑Z$�02�SߍT(�vxB�8;х�a��ð�ڀ�@ۀ�������Z��pq�"�ד⢘��<�	yȌ;h=��K���)�=����������8�O������sUʗ�C|�/����j=�_w�{u+�`�~�׀����I����	��l����u�G�c�1�Z���]*���5v�l���۴�l}ȹ=��8�"3�	E�GbI���qtp�n�`v�W� %}�����TlZ	�x撁ܷ���e^���oE%tL�W>c�J�S���n���N��v������}��y�N��{�o��2�\�+��q?ů!�~�p��N��k�*���P�E
9��:�,8���rf�sHi��vJ�l<s%1g���t�XH����-���9���Sgn ��E�/��hi�\]��nU��A������?�n=d��s�*�9�w�(�\{j
�?s@C����Oo!��� V�)�"/�n��?�k������|٬�|>+�*f0�1��i?L�������0� �|gH&C�3��{i6�koS���z^�K$�h�K�c"p*HeW�k�����'����qG�8���/�����U�0�����&��ܞ�.�Ku�k��?�4���9s��#����Ns���
{��J6l����|C�~����%�W&?�L)ǅ��� �y���d�-�g_��oW�[��}��[��Yl�v)�ڇ}� Ր���0��H�"����R�*�P#���veY�D-�o0^
���'�Q6�6�3d,�ߐ�lir�a=@��W��K|WY��C���Z���ܢ�����2@�dab��~�I�f���#5J[ve�Z�����P���ZF�I��({�Ǫ۴�
`��X8�O<�	`�Ы�0|7w[S�{��+R�o�`��=�j��N��C����5�D�T�=�
��Ҷ�G���[��� �=J�`���[�e�MUy�7��w#{&�*bH��ݼ*�N��K��$Ol�:{Wo���q���І"n"��ֵ�L�k��M���8Q+DE�]��ϲ��?H�`A�00W�x��O����;�.D�2{i��a�H����_�D�2ԯ�U�Cs��Ȱq���L��-��e�h2�?�8���<���i����?�Zz����웒�� W�~JX��8�2��s� w�a���,�E�%�^J@��Q�;\�ӷk�WE?y��E�YK�b}�Ғ|�z��$H(�O�T��?^ȭ��vh��Cdm�@���h�A��h2��A����G��\<;;
���j�cc�l�C�}D�&m�T���"�O�<Jz�ߏ���v�ܺ��O���2({0������>���!Zڀ{�-��;��o�71��nN-kZ�"��Ac�G��J%?;�"�9��]������^ ,��qޮ�*1� �à{�ڜ����;@���S��g%q;��$YH�Ԙ�V�!����uX��F��8��UЂGP�9fM~� 4e@% q���B��>�m�\ �[i�V������ś^�o"��!⤩�B/�6&��bu==u�q������"�o��F�Z���!�$�g�O,o9!?/����"C]7��U=���kW�̹2B�b��r�c��-��x{c�r�V�
�F���9u$yDy}�Ҳ��մ�������.aa�W���z��-}L��p
LPθ���z�'�ᘫ51�6;k}NH���~O4�{��[��'^px��)�n��>\n�3�����@��/i��D(�]65��o�$B��]6/��
�QR(�$�>���d̢�Q����u����Sӽ�a�E��4��]0�{���Τ��-�>�y@GjU�������@�]�Y�K�Nbg�f���ڮI�8��+��n ��zR���U��ٿ��@d�7��>�
ot��r�bG#�:���O�L팅���ȕ'BS���{c��.?����.�}��A����-4 �H�.��1�B���T~�RH�����t���E!��N��[�;�م���P�F��wAc�d��%M���s�=O�2{���\o�����A,9�Q���I �rU�;�B����i��,J_����fiJ�՝�/g�Qx���Ʊ������a�G<���?�az������x��Y�5娸�U8;�|�Դ��/7Ix�f���hFЫ���	�����] E����ϼ^���j����a܏WL���`�=�f������}s���N'��1Ԙ�h���Hݼ$����������C��9q� ��<Ā��ߛ�/��гV��DZ�}���J ��+"
�+�O�L��7�?0?L �򰀗�ӵlެ��v��t�}}���I�/��ͯS2����[�#��-"�4�x�9Iv]`wN%"�RZ�����Q��4AT8�d����i^1�H�`t<�d�����&2�[i�z��ɚ���R�9�M�[΂i1Ǎ^{H��=�=|�U�@-so@����Z|�c5�A4�>7VP.h�b},0Fi�l�+��I�r�G̼hq{Em��	M�x�D������ɐ֜���(?�ϝ�s�����J9�eQw��J�]R��H	Y�x)�䎨M¼a"��P��IX�H]��K��WR�KG6�]Xų�a&)��[�i5�Phiru�w��ZQ�A}�K 1ؽm2,#	<���R3�c�.�!��Ц�mfh���	<���oe�m�_�
kT���K�`��(	Pϒ�/�!*�I^)���ĉ�is ��9?wM}D�GV�u)y�X�Z�Ƞ��j�JFO4�T�^��Mb���O����M�9�P�{~l�r_�����ހ�N�@ `۷7C;{s0Z�?�IҰv��ə�\c����i��u����B��}����vC���FQr���H:���݆Z������w��!��w�Q�hp��>L;���.��bk}+6~!ت�p7u���s�k9���>��΅�DcW��|рg<�hZ� �J ��h���v9��[w�/a��Ƴ.v�;���`�5ty{v~@`�j�I�o�����j�vāxr�J�ʌj4�2����6mɫ|�\	.��C'��tр���=Ձ;��U��`�%ʑ�r�ڼLmp.�.�q�Ü:�X|�g�E�<�4Ep�/�ꞃc���Yl�(ƍ������$����Pa��~Ӟ_Ղ		�K�r*zy`��UyYUc�x\Sk�!{��D��\-G�?2��W��Z����b i#\	��TW����2D�KВ}g�?V̽��s�f4��BHy�:⾛���%�-S4���ToN����K�{�9iJ֡Doy��==Z��i>�-���b�nu��N�6}^�hlc�<�����
~p�LlI�`�y��Y�=���95?U���{.B>�	�.`�qصs.�6���hc��0�5hc���gv�S��_�^nVs�V�?���&��{��&[e�XQi�L'3�$�-�_6�����}�V��[�#sz� oC��!�@v�!�zR�z�)ؚեtrb�)f��]�=UQ�dk��Wf�N�|�E����5⥺x��}�߅���Q����a���%����|�7���*�Q��n��h���oU ��8b��9�� ��EM�����j�ɇ\9�$BnP*ż��<��p�7̉���9��C`L��v��RfF17s �7IJt�HFr#�e�����f��U��l�Q�ۧg4lx3�?�MU�SCVq �?��|gL�Ȣ�LL�\��z���^�DP���*�ܦn�A9m�l�-��G<�%�h8��������<m�0%��>%�����5���rSn��;��F�u{���]e2]G��ُ��񻂹A��>Lɖ`ʈ�I�Sr���n���|�,Q���.�������j��Ĳ(4L�a���x[E�}qX�?�Y�wA�>��Ii}$������+������4,޶N�jjhW����`�d ~˔��m�UO����ptM��k?�J����@��F���w���#�j�NC���D��5�t���Z�+���(�[���]��=U;DBr6��?a��x��\t�<��E�/�V`[�$�NOFR�o3��B���h8���53��jk����#�I�cu-Vx�KWp�J�Uwؼ�R��-Z�5�bLv�����k[��]EsbL,�_�E��ʬ���#�=vS	�%L��Q��ר��=]:Q���I&��!ď��?�냽Y<�I,�[�󑽆"�����D5s�D�����2F;��D�+�b|
�g���� �4�a�����Ze�*�jx1�G�,�Z����D6T)�8�i_��Z���l!��2Vm-[���t3/��İQ�G��DCφs��M�n�xW��k��T�}W�^)#���-����L�Z�+pl���9��̺U'W;�Jr���~>
�]:�9���4 U=�|�Z�ѳ���Xm���v5.Շ�=c�Cu�pP~{�5/jT��B5k�����ef㽾�G@��Lb����:���~m��)���U��W/��VvM{��hmT&7?�t��y2��T���) <.�R=]ک0M����.����M����>p>���@�r�#���'�f�\���r�"����D�EH$h��jG�x�L
�1�C�7�D����I�A�r������u��$�AڣxJ�s�ԣ��	��5~�)�+̒�&�8Up�uCeZ3��r2~#�-'������7���8'}��-�W��
c�S�8�������S��1��{���d۾�G�Qu��,��0��7�m��A~x�!pU�HW�Q�KP�i�:K�&�I�匣�,+�%_�ĥ�z��x��!�,�o�fC�#�����bG�x�}&���#�*��'�,O��"3|Y�\��6�Tq۰;#׶��$lD Ev��v�"v���������ôS��ŜB�G�:x �r��n��UҢ�h[r���j�C�������k�r��)wrZ�*撕��x8l���k������,F����ҷ�z�0����B!�
�E��薀5�����.'1��r9v�C�mI��$p�ZԞF-=��e�ۺ4�s��.
0cw��+��%���3Yۘ�$ہ _ܪ�*֚f�X���q��?���|^�I�kݻQ�&{[cwٜJ��\�U���_�GN<���L�i7��]�foD�tV0��,����e�@�<}JR7C�4�����&T��e�D&TnT=�M�9����zku�W�s$�@�m6�� *�I� �I=-�j�GX�6˭1#�+�j��hJE��A(��ol0dU������"�����];�����<��Nc] �w�Rq�W:�;_�l3/Q)h�GU<"��Đ��L|I &�Q[�J��M"�:�6��}�/����f{���3�ƒ
ֺ�=8�~^���PQ��pT(�Ec�,o�L�-M*=��H��wt�W�����?^�W��+M���l�D&�<:yZ�l�*����X��o�}�4�wzV����S�#y�h����C��D7��(8���L�uYF�¿���xv���*��N�6!��#	A��P�v���MW��c�ѯ���gr5���3 h�S�y�v���|N����"j�4H���Ȃ�<W�Ҽh|�	��vb���$�%���ݬ�7FPW=����������M�0~���A՘��f��t|��|��p�>��N��`�o� �Q�!��ſn(�߿�� u����Q۾!(�;�s���c�1���f�F��L�	9��b�0��^~���R���rXs{-��W�(�E/D����! W:�DQ�VE�G,~��U��γ�?9���/�jZ��=�e�g�����e�ˈ�pR�th�ǘ��zlOЖ�f)r�`�vU/��"+ �Ȩ��5���A۪ )�ݶx�+���N4��-M��_��a�Y�w�N�P�9��N}������:s~��-H�t�q6�u�B��M���zs�ZI���@ѴC�mQ/�0�����|+}kێ�w�d�V��Mz73FqFk9s*��܁�۱�ͮ�:?�-i]L.w��w*T�/����u*������:՜Ӭxdw'����=�&�mn�5l���cſ��%���5M1��iw�8`Y��M� �*J�
�U�3*m|U޻5u��}M[� �T�U�� pkSON�t�\�_h40�=����skR� }�_�][ �(su�t��
]�o�k��eX"�0�m�a���T����[��sѦ�v9�5����~D�>
�E�MK[�D|U�4�@�Qan}�2�z`Η�o�_�zND�f;�i�v�� X����=V�ChL�E�(�|3|���)0I��QzT�f�DM���l&:�	ᗝ8&�6�U��8\9\�q�����E$Bu�����~�};�,�͈� ?0.Zפ��f�,ק(�TVС�����}��޷����3Ts�`v��W��r����'����L��y�BN[�/�Ӗ�[3��c��(@��S/�UM��/W#蓾�d�`�"�,��f�R)C7KC�\�С�����8�WWQ�q/��iGs7�$_�]Bb�<i�G'�����Q@kNg��\x�����Z�����ӳ��nu?����B�����~�[�,X�x�O�ca����,�B��-&"�6L6�O���S����9\�����f$��̟�i��[P�@��|�9�TZ���%K��P_Q���Z^�����#��.�5��H��[3R�b,�4$���Ћzp���	R�����mFQ�^�Dj�����e�C�;c��v��psI�^Ct)�o.q�E���]��$�o��?�s�&���2Y:��*Q��(���ab�]��|�Y��vG��g�0j2�v,�����(:u(K�M6*�����Y��wلsp°�E«���!Cρ;�3TA�V�+vCH�i<�O�`��pW�S�3�1V�h���d�lj�n�6�1�<�0�jn�����Za�K/�
����/�B� ܝ_��7���Q�9�4}����
���*���ԙPr�;����e��E" �B�1(���KG����H����3� h��əy���ܛ���R�a*�zYY�9�ơ��$DJ����D�q�8(�����v�f�l"�~����"/A
�эU�%����"n�JR+h�O�Cs�s6��pofJ$6�\mP���NN�U�k4RJ�2la���)K��ܘ4���J�w�|�,��o�}�P�!��D�l:��wN7�'��@z,V�� ��l�X���@��~a��
k�Ãw!&�x�4!�9ӥ�^��-�H�Q�_$u��2��ݴȆFcT�:4 ���D���z�o�V�����9��	�5��!X�'�yw|��a�����f�F+��bmAF�5̚-4������r!�X2��	-�.b��ϒu{����M��+P:����I��~�����<.

$��q�����\{U�a��ŵ�-�s���T m�ZL!������22���� #)���[�e��u������	�&{ ��n���l&F��b�L�>F)�w�4�o�:��j� �Hb�;))�3���f��Ƃ5�Ž���9 (�Lߧ�>���4)�ݳR�P�/�^mv��I�w��J7�P�#��D����e�Wȱ^@S�混k(�GU�ĮY���: 15����Q-��uC��˸gu�L����Ė�eh4��:��[���)yTM�H�1s�J�nX�-Ö[��	�}��\+�?�$<D3u�n�au9����0�C�5�r���j��-. W��[�>(�����ꟛ�9v�^6,@?Q8_����_u��x��/���"����oMn��� ��Nו�ȞX��X�&1�AD�2��������4㦦$8�+���10U�U�\<ύ��ZN��B��@�3�u0��1���8<pN��5p|�*1/����M�-�%$��ں� 2ۉ�2��d��6و��P�/FA9� p��*��cm�XM�ـ2#(狻�!�Y*R�9��Vű��e�:*CVf��I�`��wL�� Wk���
Y�mAs�H腪����:�x�]�C�P8_if�U�2��:ۍ���,�Rz���i�`FO��k�j��MI߷��G�[�q�a_���ʉɺy�ЈO��j$�~�tbD� ���4����Olù��R�0��Q�Ձ�Q��jhA�T�Ak�X=4�LfD8R�:8�a��U���y���X�`347�c����YN��`v�X��@H=���!<N�o[B���>���6$���gz�bV�oQ�U�	B��k�0��*O]pKW�rŔ�r��tn�'����3�t;�&ڭ��d��X��h�P?ɖϖ?��}׳mԟ"Q�d҄���g����$?�D� �J��k��w�H�^��/�Z�8D�{>2{^�zz� F���D�x�[�w�)�������t���c��b�'H�eL�,��&���qyv��6k��&|�^�Q�T}��΂/\9����29�:�]�"����yr�/8G��	�q7t��f�-��վr�gA[_�����j��y���Y�ܰ?�@�ρ��4��e��cй��Ĩ�)������|��	����?�QѺ9+5<�d+�� G'L#^�#%�e��A��``�\Z�6ț^,�CL?�<#mKB�RŴ46�8�Tz	�1��8ɐ;�7wl��%�BxYߩ�.���t(e:��P_�e{�]0��A��z�	2���-�怔[L�8�[�/�"V�=�?)T��6�m�X5�KFe �ؒ/��')����<:�
ɼ�g�9 ��.��_���!�$��+���b4���␚^E|��yP37M�U���l` JH����t�'+���].���jk.�Ŷ���O���r�#<�|��²�zs�dߋy���!�K��
����������_Sj�] ���;����1h�j��m��,}�OS��D?�g����m�;ډ�\�������i\�^J-���6���n�$ ��{���Z1'u'�!ʇڱ$����u�?�� ��iɑ�N���cO�*}NAvɏu	�۞v�k ������ҽ�G۠�j���E�����]-�j��-��u�.���V��v��i�����L�t�	�� j���6�W��C��)�@3.P��z�-J�I�������F��2���<�K�������S��M5f���^��h����&�C���E`�k��ӂ�Ҽ�ٶb+���aW��_/p	������aRP���w�@�N���I��/|y����
�3%���&V?����`��]d��n�S ?_IrcphW4���菣t�ְ�*�kԔY{>&�j�ԯ2������w��B����4��f�5�r����`M8�C��/~/�q�ʅ��<��M�<ߨ�l�~�T���^J�f+ ��[*2_Z����ۘ�U3
���B����چ��|1-��RF[�:�z$^���C:��O2��>�L}�K^�8��{{����k�2��^�W�����wEu��<�XVFɯ߳>��;�
]C!��ߙ�:��,�MG=2�~����?�9c$��L�i�d�$`���:0K%e�s��n˸���X�J�o�׾�,�|�	�i*��ky[Ԫ��;�2����c���	����V6E�gw$J���F�@��|���n9�lK��f/�!\���Jnk}L>��U�nX��>外�$]d��5�l�P�^��&#iI<�khΧK�R�)�pe���K���?�C��h<i��I�?Fj�ɪ_�f�4�!1Ty	p̐/�uf �F��ais�qD����ϥ��kg�����Bl�����)�{�yPU��<zy��Q�n��u��>�����nH�c��{x�z-����Ҹ�b8 ���$i .���j��E��z\ڦO�$�>2C�ջb�o�p������ž����}�2&�L� �o:�{� �'�^��ƒBIS�����ط�Ak{���z?��`�r��l���iGA\���^X�}p�B<{b{��i�HZ�=yvB��ҸK�k�'��j�%O	p/�S66�Fy�.��x5�M��B�;�����$��1��w���ϴ��mI�i�U"�6X7	�}3#�[�5���O��� ��ٚ� n�,s�����.�_d����;-,��ڦ����>ԵI��h#�9�ܩ`�Ź�X���ݼ����^Oj6�OL����ى=V�o!�����XzϜy�r�YD:HG����ky�`p� 2� �o�L �cy���9�� w��y�8RU�(9��a�m@3�P�yYe�,��Vs���7b����[RaS�hCߤ_�|��TqXeӾ�r�1�����G�9�C��8��%�6Y�W���"��p:�w�����Q�s����{F�;��`kxΛN�ʤU�����	Ls@t.�M$�pl9)n1u�\��O���{����:"��g�����!a1D��Җ6�Y��/X�6>:���p�q=���6����_-�Ӕ1�b���e?�r�m:��Xd��S�6�Ȟ�2��8$)�X���6٪�Y�j�EK״u���[��8��úL�L�_R삷oĤ1@������}ao.�tF���Vۇk^:�E<ZRNw[��nh�a�3�w`�i������kE�;��%�4��#Ve�8�Es�DI9�;u�2����2ɳÂ�x�֣�L�
&w]Y���w�I���:@ƹ�\�{�Z`������+��$�0N�I�{�t�bb{j�y���Q��U'7Pu��������7O�a�S��i`d�]�أ�cw�����v�O��M?�O��[��[|�~p�u��;���U]����6soǫ�s�,7�'�����*�9˦=���%=��� )�hW5z�&3�`�� T������x\�i���L�:az��d���E���T%D�||���m��.x��S^`�݊|�IfDkT��[|��f���/ڷ4@�Ђ+�,��l>���P#"#�d|�P���9	�Q�Y,>xf��*��o	����ԧ���_?U�܃�gݦ����ܟ<{V	�R�b�U�ܳ�g�����y�
�N�@ȏ�oW���R 4g��>�h7��NF_'�\�ԊFj�-�����L�daY7�z'[�����2iyQ���}a�e�'�4�Ț̡����2$�B��J,#������D�P,m��UNmIxj�#F\�^J�㫣��75��y��֛�Y]*����Z��O��zJ��{5st�q4�%m����I���+�����Y�d&��EH>�*��x3JMx�yE��آa`
�ݝH]ؼv�{�y��8[��C����<v��8^vɥv{e���7��ش�����*U�����w_�Y�q�m
x�:y�x�Da��B_CI�'��E
���1��0�Vc�Ǹ~��5�U�t��*:UCl�%D�T�T6Ila����G7#���7U�������[R��Z�r��n���g���4y�5��b��y�w�����R����K�Z�H�bfW�NeqH�®c�9��^/!�̅����k��+��f7^��	E�g"S��kΉ�Yyc���u�2��̄koV�FƩ��Zzg��$<3�ڍ0u��;��a��Q|ݗ[�^�
����<e
<���.��e	QT
��rֹ\��`��+ݍ�� I�Y� ��m辈c�Zr	G@��H��5����Bxt������������yq"����%��[��/V�x	�)#��('��^t�<����;�$c΢� �qyuQ�&��U�{g)ih����Z@o�3�[�KnH���w\`���sՁGJ6@�c��`@�ᢓ���"�nV�}�9 vd�&��#�1�QV��2���=�!��	��T�ÄS����q*�D+���3^d���NnP}�W�?�-�ߗ~v
��y���քnf���s~�V���ҭR��t+.)�3G� ���t�!���ĜK��@�[1�\'���u���(%���Qx��R�ɽ��Td�A����i�|_��#X��c�F��*x08�.��d�s4:�J�꠰��b@�(%�[<4!WVZ���x�:	==��)���vȩ[+���l���ի)�Je�΍���.����4��Sr\B�3K9��J��x]����NL����iO��5�F��U�~b*6_��9�4���t�S�����V�	v�6!$���b�@Bρ���+P�ͅ�.�ܺ�G�S>���)Z�~P����V?U%��NUA�u�M�BuI��6h}ËX������+��Ld���w%f�'߶3m�| /�y� ����X�hPdV�E��PAr,*�Z&�e	a`鯮T��}���l By�1Pl6��as��rU�(�e��H��q�T�_���_�2B)�*��ё� �)Z�������d���:��V��#�Lh���%�a�)rD����S�ˏ�����O�mrs���a�������`{1]`��A(2��7OT��8[�s�d��ʏ3mgQGcZW�26�YFߢy�pհ��'m옰����-�l�v���6����0��E�ެ�7Hgx��$�ee��;*�G�������}��U���
�L��-��'�Wx���t�扽� [��|I���;�Q[WUX�����0w4�P�==qm�?:?�K�p�DS[��_�[�~��!��(��1w�.�-~=�7���yѵlp~y�)��`9���1_���c��%Gv�(��%!X#e@&��M�����5*�ȫ��Sn3���E'����0�_B'���_���ǹ��8Ķ�ٿ�/eYC�%!kt�s��ύ����xR��W��Jϭ?��$:?��K[�[K��&����㡒���2�k�:�"M4.��?D��p���M��f;~䞾�k��_Erԙ�]o�N�p�q��B7yp#�@Cߗ���E*}|6?-?v�,c|V��·�A-B'�\X�	�A���TE��0?�����F�$�h���ṅ[a����h�6��ɔ?���V�zAUo1�P���� Hx��v	���,��U��^@�DA	$ζf[TP������
j�OWڞ$ dprZ�4:q]Q��RK����A��K�&�N��~�R�r,�����<
����W�tk��Qu7]�Q^	��Y����>R?Ϡl�\�X��N��|�
��{{���gů��S��<!�7>����) =W"�YA+E��yl/���B>�1~s�!ѣ~��5��7���7��(v���R���	�bG�J`����*t�ȱ���uq��N/�Ʒ�}��Y���x-�FH37:,t �#ʲ���ںDGo��� ˀ��Г���2�)��ǧ-�zV����3����GXՏf�!�EV�xb�����6<���6ZL��ψM�+�%s��n�J��<L*�V�T�$w�!�cUL�y$�/%�]��fU�Qp(��`�)T#9��P�q�o 3]P5nj� �*?�uHW��'~��&��}�փ��$�a:�,��W�D\2=�����E����ֻ���y���M�ho��riEj���4թ ����#�"�Œ����@�h��v���G�hGu���]���6����Z!/��O��>WQr�ܯ3�����_S p}P�ԨB}ܽ�7��r���!Me�h�9&��v~�e��k{ks�Qʁ�+�}�ՏF�t1�"�q�������Fr�s��U�"ϼ��zj8@��)�N�H�%���{Dn�Ӫ7e���K�T���k\5Y�+�;����_�3����v�s�og�f����V�`ѫi�[���0H�\d������ �Nt�T�% ���d��6xU�FD�j���u���-5��	�q�G�Z�h�DLڬ���p7��{�<�nP�o�(�Z����]��b��
�~�q���dc�ٗ�|�B҉�|��?cv�,���R;a���6�� �1�<@���q ��1U�������S�}x���
�UPm�E����)i�}~�ON+�N�#% C�~y�ysF��+����0�_=z��}Q����wψ��d�O�q��J�G��9��F����!��i[�|�l1��l|W�ܜy�7�/[ѠƜ����d�����r#(�ν�_�����-R�f)�<w��d�[[�=��<����[׳�6�:��9�Б$�j�Zț���.v��1ު��������*N;r�&Cސ��dC:��]��T��g[?�yub�z���c!��
&G�N�~|��;���Q_P�-k�	CD�OU���FR�1~�E���#�-�����2�� ຅�܉H�� �Ff����U�������[�儁iO����C�b���YwM��NhûƏG�@��&����9�^?.�ł}C}�a�)�i	f�4����"�R�e�7&� ���c��6*�B���D��������f^>6��G�}���:������r��D���m���}v�{�&p�����A�E�����XQ��wԍ�:��h�x���Ut9�w��Y�EnbY��(J���;��'�k9�H�uln����Vk*�������u��h�f��Q��ֿ�.�p�c��h%X�v�M���ü�7캔K��x�i�P��R͗��x�0��F�{�C@Q��.�����_��6	���\X/�$�b�6#)�1�B�[6���h�o�?�ڙ���Ğ՝�N��r��#!�q�n�^�U��;g s0Q�p*��/�ϡb�	A��a-z�7>�k���mۡ� (�z��Uߵ����0��f._h����k-�� I(�� �����*�7jҭ��a-
���*����P\���,��3aZ����r�#19�÷O�bs�1�*�$^A������ԭ�&�M}'�%m7��ӥe~�^(�u�ёW<zO�n��@ݙc�i�(��0��'!�)��bn�w���"_G��K�G�3���t`yT�Z�ę	����,"d-��VZ��'�(_��b"+bl�'�A^�f�)�nE��ҽ
�iO�S�zZ�H�O~&e��#LG����gA��k�Z�ǩ��)�_����ΤG�����%R:
T�8�#(=`�2�A���H����� ���`ȥ���\� �J�y����1?a����G/�ԅCqZb8d~�'Z�[4�0�ɜOh@L�@�1��hH�Ν��Ɋ��\����J�}�y�K�Y2����.���:��}Ar�����DA�������	��#@����y��j������g�����nz�s2Ƿ��n-�{9�*Kn�(�{jDGfwZ�U2�h�t�F6�Ok"z]��&�.o%Au˿;j]63���#���)8�0��HV��@�B �Ql*��*���F�qCBp8QR���2\4U���aH�,����z��GeN��E;�ׄ����U�f�T�J	�
?�#��8��Sd˵�Ƈ6�=���СG18F5�[b	�=�z&	ϓ7c�����2��\��iyI?��z4�3����b�w�c� ����'��A)�GT�EM �����ɴ-]>8N��?���&8�pڡ�L�I_���ɴ�����ve����F)-R�Ċ�@y���7.P��j��wTx~�L��%��6vG�@�n���@Fy��L��"�w�t�)EG��T>`,����1���Dt����c�n,Fm]ϻX4ز��^F���|���Ԁ3m����uk^�V�tb=L��k���|��i�Aȷ؍1 Tw���V��A��q,t�/�T�-����)ʜ���e-�G�RC�k�33F �r�K���AR#^�ݘ�����_�'����Ju95��Wv�����F�-?�F�S
Ed��)SrW�Z|EʉM��(A�݅�G��(%U,��F6��f[�rt��[,[P����fԎ��0ʪ8[�C-1��F��)0�j�	˰�]1r�z��ˠ����r6���=v�+V3'�O�,�]�r5aEr��ϦG;��^pF�����yA9�6��v$Թ
�֨�Q��2��v�M"���d�2뮀(�z@���߁�m�lxN�*�nNՅГ����Jq��B@1oR������w\V���g�[M�rW��-�@��`�gW)`��8$���,Q*1� ���t��0���s��uoo��^��)���Z\����G�x����f5�p`�?գ��W�w^��E���#ofF�`T�?��]5�I@F4���~���;�#�x;)ɜ�>��`iY�\���	��p���Ǟ���$`�GDm�/�QxbV={��̖�Ք��ͫ������	<���H�s$g�r)Z�tzLݞ/��p��é⛊ sM	��yo�ԑ� �T�朷��/���z���t��Y���![�2$��1<~�]
q�b�u˒�۷	�a�m�B���b[\���˰�)��	z)��dt�)Pčo���Ð��w8Q�g�ੀA9" %�t����j�������h7�ϰ����.�3H��~�R.q7�a��[r|$�Qj�y�$8�aw��И��xzl7[zM���g�֔,���������NH��GI����4G��^�-����Q_8�,�k�i��/���e`����J�����D����s��m�º�ⲋH#=T	�L����oOV)�1�+���om� E$SҢwL"���>��N�Kf�����j�t�Ĩl��-w��;3��>�A*�wX���~�2+ƩI�V����g��aˣ���DȠ�}s����j	���$�i�y?�M�&�u��ӆR��Mp�2����
�>@eY>�w\�KJT�*�$��F��+����y:5�xb�G�2��{K�w��[������(뻗�<�]��#'�&�H�6���R��+���9��Nm,;�SW���K�`���7�[Ώ��'Y(�h��q��)����}�_�w�@�S'�n~a�Q��&/�Y! �5��+��#	�"��;2T�'���SI,�<:�Q*ޱ�M�.��*N��h� �^���c�&s�u,�e�k�2��#[#�CL��q��)����O�NP��sg�:���Hl��ȁj��큖��0�Uϲ�P�04X��,��o	�Z!��u��@Y_6^;�r���� ���%��R��ݮ�X��0"�u�&SЛ���b��rd)�Ɨ�6��&�Y�[�j��-%U�~��V��<��ѕ�MA-#)$m\�t�-�SO2j����_��ջ!cU��z�ڡ~��ה��I�/?Q�u��]6��
/Q�i��C�T���l����QV��(r0�J/�k�.�<�"K�KR�N4��v$§M7x�y�zS�C 
tNK��w�Z�0�W��(��f����a�T>,M�!j9v�����N]4�Ln(Ӂ��f��^����w�ɴ>i1
J#aq�7�rЭ���u����֞��04ص�R����.�m7��>����u���[���%��>'��f,���'�)o��jD�^[��z�ś���r����ʻi�����P��?�H$(Ӂn��4e��������b�n@=�'3�K�r9������H4�'N�E���N��p��z"�B�Y��ⰈyxB�� LdX�v6�_����]�vD%מD�<JM�8�Ɋ	B7g7����"��g�\��%N��� 0��b[�߀|�(�B��EWu5aEP| �M�g�y���zc�lS�.�~8&	*�>Y������q%�e�F�%$�I��	a�IZ/$�v�ȁ�����Tɤ��;�)@<2WF���9?���>�� G�@�t��)'&I��Pr@{Z1Z�β�/��h����>xr�?�(�-{��j�8�nq�`��+�Hq��>�ڙ���֯l~tiB�eŝp�3����9��XP$ӊ#H(��7�}-�_V���2����t��_ϮE�J�1���v�H9��+��/{i�mf��Aϳ����D��h�q�F���@���C���~Y�bE��\���i8�TK!(����G����U5�=�^CV鵠`�毂8�)lú��Db�v��9\�|!,Q\fn��d�fo�ײ<�WM~5�K��3���AG|���f[���	�f!
-�	E�h�Iu�NCz�j�R��:�1C�%;�	.����G����0�ZYރ;Q��3[���1�Q�<�A���:��e+���.Ŗ��4]��H*`����BGy�X�`��� H��Nm�g�ۆ��iG�9٧�T�"��M|!�����ʚ��)�(dF}�w�?ؙ޸��H�X^|�����`���x�nFq�6�e`P�V�.�5ȟK�[��y>]S��W'}�wt��V���6^#`g��JBg�&r<.S��ˌ��s��x�j���S^�ɔ��k8�����05�'A�A��3���D7Ͻ�ޚMKk-�+���W�@9nX�����Zz�/��$�j�-Êª�f��Dp���*ȃw8�ƣ1�H�Gk��0N�N���9���.��~�$J%l���$?�Y-�e���=0d���&w��e��5��cn����vc�:$%�G[�>P�l��˅�&�E��濏I-[�M����v:�x�f��g�z�=_�2�[۟TB�3��n����!�� �Gl� t�tA+bevp>w:*YU���hJ�>��@=��G�B�t�\��(v���И�$�h����F?n�d1�U=$�?a���W�� J��'ߐk!���ً����b)cw,�w6��{��`Q�c��T��\DoJVO]�@�bZcE�m�~a�Ҏ-���k�s!�ГX͇{=(���&p50�b�}�%ļ�}P���!G�/g�^��A�U�3��{d&�R
���-�z���œC�m����YM¬(��̛����A�ċ-�Q<_�����
#ko" y�{~�a槟n&r��"�O*��3�
w)5��7/�����x�c@��ڽ��K�C����$�'�K�z��
J(���F�S�����Ù����IT����[V���
� �$[ΰ:�"��%!6�}�`� @
��ܲ71�xk��ц\�w��>�_tg����$$��B~8r���ډ�`*kޑ�υ�I�iW�6bn�������9�{����Q?P��.D^��n���`+�BD�J�!Ҷ�΀^[��NW.�ban�o��tm�tq7�R�4/o�����?P��'';�=��_|�Z�Rb�ڸ���5����)m��N���܏�y࠘�]����;��kaW5ǆ�U�f�d�U'y�{����>�|�y�ÃKtN0��糂�nU�_���g����>��0��[�V���v��-Ēm0}*�ϥ�^܆e�n�JlL��X*K��F�Z5��*m��C*,��ե�~�f#Iaў�cR��YW�������ס�v^��Z:U���y�3��aG�2���!=K��>q����꼞�ž�IFԟ_aԳ�NM�Ǹ�^Ǽ��9���4���)�T"�P�v���,�}ܾdf��n�}��3����ntXo�!� �VYgwj�R������<ZVz_$����J0|aY-�췲�Է���&����R�lhj\6��r��	υ}*�p5���Y|Qb���C����_\*^���E��ܖEM��H@c0W��L�䖪lB��ͥ��ji̿�ù̽��&`gg���j����z�x�%I���\��?���X
t�mϸV�>�!��D��эV�`7x�
](̰��*{-J�"B��͖_%���F��ٚ㉞`��{��]�p������_�>@�ž\Rn�6���a���R���YjQ���a�V����]�9�Ş�mupxԛ�jf�$��9जO��ֿl�+r@���m�rw��9`�BXf�1���wcKr����H��=�X���j�_�9`�L��Z�Gn��ۿ��-�}�����G2\ǃ����S����+t�$O��ŗ7�o���DH�"o�&m��̑���&��>�jDɄ,�TY}��
��G�8��}��@ʍ�q,���@ѷ	'����@�C-����:|��i7_E��K�|1�Q�����?$~�4g�4{�c�wq�'L|"G�9!�r"�0���'�-:BG����t4�#Y��)2��[��N�4�!h�~�Z�PF,��K�/ ������k%��~�gK���ؤmkC��VF�t�r[��U}�Jd��>Jřde3ghMn���:~)�^��m"���f#OG��W3,���b�-�,�u�d̴��lH���+? �

��Eh�t��3���u�Pv��L` `,A�!X��Y�ԇSU�(
)T���.�c5Ɯ���r[��B��t���B!�+�d�r�yBx��S�RW����7�}�Xk�f���'{S��`��\�S�p��ܟ�G	\�K������A�>rc�k����)�z�wgT)~�O�c��怃���x�2���
�J��KI-߂�2LE�\��/|U=���6/���@�';@�:�D� ��N��3���|6�E5�����*T��0�Br�Sm��P���%H}�6XI�DL���v�b�J~��g�FᲵ�Id2�&�%GI;��Q=q �G�(O��gAC䒰��0��`��P>U�d�uz���U���b�>��ķ¶	ϐ1l�8����V/k����8��җ;�.8�/M�t�;4|^�7P�?���)�b��V� �?S&��<��K�(+��P�;�4�#���6Y��
a^0�\�B�f
��k�>�LZ�;@���S��:�_���i�N���P��0{��-�<ۼ�Y��"C��Vi��G�2����s�u�DWSPG�:����ݥ���9���I�
uF吏�}�U��ؐy����S�ܱ���E��Ӟ�x��t�شU��v�1y�E(��eߺ	  �@
���/�t�ߨ�"P�h=��5
��9x�%��T�%�bA����EZ��b�c��QU[Šv���iGb�H�qU��)��2S�Ϙn8r~�?��Dgڇ|�y�f� Ӆpݸd�>�SuB���{��$	�K1[F�GB���r�p�׋��i���}��:8��٦,0ixL����=��b��|D9�Q����m�Z������_4���h��L�o�ů<6�
�
P�t��mv����Ε����w��e��� �cWM���pg�#?�4��Yri/�1yL��2�T����v��W:D�ȹ,������E�բ[m�������>? 2U�A���)R�A������/ew9�%Ekf��Z��	�4�p/�gb?���Ӫ�&`����Vn�)��{�s
 ��b?L��@�φ���j��z>��m:�k)��WD�O���L�5a~p�Kl���� �f�O����5B/Zy�)�DQ	��ǀ�H���0lbk��-����Ф��9�'�V�Վ$$w�?m7�L���ƻ�gm�W.�r	��2�
�"�����?����po[��#]�R��y�I���*�+�d|W���ŉ�G��G?��í�<RnX=�~.�o�X� !�Vu؏y�K�0>�j�����w��a����uq���y�1*O�ʀ�|b�E/��x[)!k/��>��萎� o�eƲ-T��[�>v��"tY�tP���R�uq>�$9;�AF�+b]G��WT�e��l�����`%��f݌���Q�(;P)L�IН/��)�}�: ��?ğ:��D�����4�EƘ�i�o�����@��ZQY������9�+Ͽ2�>����D;�/,��-cGa%�d!��S��6RR@¾����(fhZ��zi�I�Y��=�o�:�n�N�t(�3   lH?�3l�Tʼ�9h���Qz�ʀ�v���5�ٜJq+�2�R�$/�G�E�2MZA2GB����8Z����ݞi%G��.`mߌ�#�o��K1C��{5���������e�e�6Л&#%{-Q����'f�A{|	�@I��Ԯ��a
d�\
�v��-!�����;,j C�>�Ӿ��]�z�W���⛗ɹ3�!dST�9��X���ĕ���Ng�w+��U�S�B���U=���p�Xf�{,���(�TQ�>��>�#����BYĶ#�$LH%bP�����P��(�?e��@�èȰFϤyo*�����k�v�`>F<��Xg���nOXQ���-\����ͤ}�l/^�̙C$��l ��娇H�(�DޙU�m	ÚFɐ�#e�a|���Ld�B�:�}z]}�\�uGHM'Z�����xM�G���UR�T�/E����˿E!��ؽ�Ѿ-�e�!���������u��bhW�_����'�G!�_ى���V���h���B����9�t)��Z*���۴��R��x������Ft�|�8��/IjR�B���J�L����m��򺾼F��hS��#�]|�*=vȂK�űr�"����x����4ϐߦ���5n�iׯ�.4��'3�$�)"�s̕e_b�.;��uB�T�c���̆
(/�q鏄�Dʅ�K`�]���Vh5Gr��&H��UY�����4��v��	yrȟe��w���h�@6��@K� )����ď�^�p�ST�M�Kr��0���	[����Ѱ�e'��_��}���zŧ ��]�F��Ut���֤"u38,��݃n_N�Y%�Y�܂��Gj�_MklJ�.����j4A�I�[#ߟ����Jܫ�<E�w˒��,=�� �`�X�*fJ�a�M���-�%�SD˸�A)���q�[�F\WY�khRW����,P�����!�Z���ݙ�y��>��bP�c��ޛEf����h��#�E�7!��C����u$f�6�K��ܜk^v��<_��//�k�΍]�&$�k`s�m�֜�:+,Z�L����(F0�Z!�F<wz��%����sH�Od����O,D9��V!~(����׆i��Fշ憝VK�c�I��#��,0.� �/�2�e�М�t�X������� Jʦwܻ>ǫ��B����h��n�8Y7�N}mo<��Nthޗ^yuÇ��ن&���gC��@0�lbJGԱ~v��?���u�6�{F�BШ�},�؉��aB�s-\�z�u����b�Z�7*'�����6�ܚf��G�G���
r��{���m@(Mv�֮A3�(�$����A�W,��[Җ:b�9л��!����U����@F����@,yp��^΋��n�)��U���W��h�.��5�8ſmt��`]k�G�WAб��q��5���t��ʐ�f� Q�;/=�H2ic̪�gr �`�t&����Z�@\r�ћ���TM� ������t�%Ҷ��$ȁ!�Pg'1��Npz-�Y!@�P��<V?�I�:���jRNP��)�|HP��E �){�u�0����a��X�&T�ޡwjfmc$�&����(� ��+a�ث�_������k�[L��t��w�}v�+�fDc:\����}ʛj�
c3���L7�f|��x����ʮ�bY����n(^�u��#ɅP��E�x_��=�@y��<VcR�v�w̵=]9�Y�u��{�$-�5w�}�`nf�r����k���8��z*N�a���-����TO��2&�Is�4��W޸~Aж���N��c��E6��@.�̧c�����	S/�-��F�<۸w��?���W1�����S��n��cRņ����Be���F���qf�s�e��g���ׅ�3�L+�0�Qw�Y�(���5�g5��`����9K8ڼ��U�)pG�9G}Fk�s�U?���w
��Fj	0��Z*8��sӷs+���p9�63J�QB�>��1�+^x�C�B
�7��æ�<.�����)�Z%#��Q1���n܄�eq;���f�Ň����;T��j<@�oNJ��V!a��Cթ���M`�5q�w*�г��id��� �H\�K䄢S�i���l��x3�\�4�}偰����jP�&D_���r�8uv5C�� �-�pa�?n�p+�J^C����$F�/ɺ��C�?B<��C�-�Ȇu�.PrsM7ؙ�Xi��վ�]S-��"I;p���'LTSP��Qo�׍jY`.���4��@B��:O���B�aJ�����hs�@���ɮ��S]�Q{XS�(�vO'$�U��);�^�vi:��S0n ��\��)in�ĕA����f�M�Eo��Mb�H�&3�0E^��T���̓��񳑮.�����>��y�@�l���7i��=MR�Y��p��L�?�_�MX�J�ꀕ��;zq�֤�(w���lN(�Z�~�Y�j?4ˀ7��R�#>��_R~ou�Â,��[[��;�3�1�k���_��1�~��� ��^,�$s)��92��T�F��Zy�����~VB���1jEKj4����F ���SoH�qB[�`�Y_�g�Z������)�,r?�����<����A�W-����Iˋ��E�O�2P�܂����' ��d�A���K���R��(�pZ�wVj�0n>34__���ޭ�q��ːUMl���*h�;{R����cZ�&;X��G����$�5��~�����kR%�ÄT���	 ��:�~+Q8\�v�q�����/��+�\X��?ۡ�'��LO>�� �Ҍ�a�n�����-P:�R#�M��Q&��b"�<����#��K���Zw��e_f!e2%����(<�����w�i<]^u��v��z_VE�O' ���R��e&}�a�ܥ�3�������	��M��XR���������4�CK/!��#K}V,��߾�F{����m�֩cʰ0q��]CH�&-e����ӯ/�aC�%]���f1@h�4D��e�+c	�	A�M�*y�T?��dĀj��W�@�;I�E�7����HNb�ĚO@������؀"5d�v��R*5�/�^�E�PƓ��U-��2��L@��7��v�I�2�V�/�>���̐폃�J�PEfE�(��]B��	��u^�to���wF	a�-Imq&�* ���ؘI_`��),��Q8@ӄ�`�HNq�*�bs_n�%n��|<�S��~n����'�xGFY�z����
�bd�g)Z�w�£��	�&��C�!]dz5BiZ�m�4���Z��#i �|��3TޣM��itT2�u��x�F��w>H�����]�(i?9��+79o��O0@ƹ��`0]u�VB�*PƊ�&�+)^�V�ۃi/��aK�� W��?h� w��q��U���K��ؙ|r��n�Kl;;�ҝ����Έ�����%����a	 ��p�,����EP�K~deU�:?����nג��܇%3�е���9@a��P|;^�߅��TG�^	��_U}��!Н*�)Ę�u��I��Ef�HU�փX/���v7i���f8�J��LG*p�4Z�%C�C�p���h�`Q)�b�|��l��R	nuG\��t��5*zIcT�]�t��_q��'V�݅�}�ڜ�4��r���<��LF���Z�=0c�Rhh������Ɏ0�뼌m-�3/���<jNJ.�c]��8i�"�5����v�cP:��nV��O]�#�S���Ƶ��;�\�S��+ �M�9q��-����56@�\���ć�n�2NR���J,~4�������_�jI�vw3=,&�;��!I�Ưs�p�չMX�~`P���UL�g�CȮ�^ؙ'>�*��J�����Mo���֣����	�+����%�t4�I7���E���]��'�����Pnf'\ǆ�*��Xj���Y��w(��*�
OW�����u�B/�����aG��QRj�
m���7k ��<:�ũB�W���4��^&�B
"�Q���n}�Z��8<�>+�ہ�
~���)��C����s>�}�7Ҷ�ˉ��1m���5��u��#�0ȑ�7�
Yo3>�P�r�M�I�?-Գ�c @>�<5�a{�?a�۔�-�>���S�32���)&=Q��ঞ�^�L�3����xW��m���3IPI�}��79 ͬ4�� |{���`)m�_�I|i*���jA�nI�8Xp yV��G۶/Q\�I��[*5�z4�%?h����S$�3c������؊u2]Z�Gx@oi�O6�C�¸'\�^�@cUƯ��/��>Ãɔ���1? ��R<�#L�({���#�EY����߆����M��d��|��x�7xk�t/Pʎki�WO%m��P	{al2���l"�nh����1�a%'�I��KZ�����zF�h�@U��P�M̎C�{0�jϾ�ᮮ^���E[�gz��M�C�e�4���7���Cf=H�F@�����j��g.�XY��ߓ�㞭I�T��,�,\m0Z�I���:��Q�r]�@�w8358��SB�<�Bq�3fK6�G uI�b�d%pa/t�8I���VH�u�5Sj����Y���"{��������&��� ������ۘ,��?|֔�l�Eҙl㥌�Z�<�,��:q���a;�t��^^~�l�$�Ug��!�:>�z�
T�5]�zG@������1�&b��s;?��K�g�Lc��1!���Ч��eT0x9~s��dG��2�v�u���8�]�L�{���*��R�~�F�n:��I陠�IY(~�aB���M�χ(U�n�s<�;�! n�;�qvކ���x�ݭKF�xF1ek�w�#��&C�ڥ�kU��%�
E2Nm��/^?��OQ\`BS@��7)���~�י�NR"�X�*\�>��Н"P��k���m�6���o����f�q���Z��Et��]���	?ei��J5C�8�b� T�@�r���m��L���~�x&W-�i�Ѯ����|���M���Hj i�J�N�D�]�9$��Bv� ���mY�OW�2^o��L�Jj�� �7C�p	��z�!�q�FΦ6�|���
��)���c�]k���FU/ם��m�_@Lk\�L�T�C�Or���-�i��BY�����R�x�e,�@d�2Ii��a��ue8T�s+�n�"��|��	�wg=z���$V���D;%HT����~�� �0�1��(��}�]�.��j_֎d�$@�C�ٲ�����h����vʩ�`
��ŷ����̧ �C.E��q>1�nuX�����nT��#�V����D�9b�&m�U�"L��@��ȴ#)#�	�$����3Kw���8��K�Ѥ�t�J�4}_�l��0{�qf�e�v�0}���;:��wH�m�Z�C���~�0���|+r�� ù��?X`۹����U�m�|��8�j�<C_����u��M�␏�����X��n4ǩT�_�ހ��dұ��<d�/�>r�h���Z��W�ͭ�ګ��R��ߔ�U"�W.ݔ=c��'O@��zƸ�I�t��S�'�:��^��WjV������Y:BE��1�r!�Ky/�uրP?��8�svU��y�U'�*��I��PF�,g\D/\���%%)x��3-U�1@G�g��ض��ZS]���BT6����2�k 4�Øܧl}W��\�hRMPڥ��{ ��۟]���2�x[W��n��������G�z��M�w��A�[������	߻y����Zk�Zdd�]��ʌ�&��R��O��[�4�I:���}M�bؼ���ף[=3�I��O����	�abH�L:�����,w�y9`��hG������4�p	+�sh~���|��N��[�7����c~	� $n/~_�k�>W��V��?��7��DjַRãsq���m�y�P��P�����-��i��a�ڱF5�ґ"�
^w�H�*��^�ք��p�rh!9�,=/�'�mv�u���vO���*�]0�u�aW�۝M4HTP5{������.��>y�����X�7>�6�\|�{Bz�h8��	�s5Z�Mq�Oi�b�2�Kf=|�A�����t��o�e��j��`w�C{-MW��Sg�ݸ�/#��r��`)Ϳh�����:.z�\iW�Z�MJ˨��3�_�5Dr�G9UI0h�s]*��T&�p"{\�E��%9�Q��D��Ya��ɐ��L���%y�|���+<�-m?<\�Y2&̬ S�u�H��;gB,k�Ĉ�B$���\5�4�o��:`�濏h���%�'48_�r��0��-�gP�T�gV4�MxъK�b��L�I���D��1�6q#_�md�VI;X<Mő�~��`�0~�Q䀁�!�xc��F`�sV>=��%��L_R��Jm�&�]�_ �5�3 �%�t�5s�4�%��y���s ���CT����%Do�Z�,SP�U.	�)�ҁ��ǀP��ߓ4������ԁ�I���CT"�T���P�>�ff&��ċ����̺I4��c�В5��R �� �X�u|?P��cs�Q������Z �Z��������
�@߭P\h����Ĳ��2+�o���q�ο�R���\ H�㴕1;2���Q�&�`�V<��������x��T�L�8c�#5������d�)Y���UÚ��U7�8�	H���&LB;���b�*�����a��icz1������y������|3�[)��&�ϧ�.�1�)~�	8׬��7�g0 ��mE?fs�5m�n�z�|h��C��;6B��\�������.z���E�:@�
@P��j��D��n;x��6����0.��Yj��5�@�p��{���W��>R	���u�����3�Koߛ��w�~?H �#�������H���`�|�����}t�V�L�L�V��=a�����v�ɦ���
�W�*#�&��"�rF���|R~���q�k����^S�����ZwB秠�� t��N6xQ?)כ�Q�G��1�H���P��'=�X��"LZ�?�-xJ�<�+�k�:I�Oa_��e=�+���D��MzVL>����oZ��qpr��`�.Wa���2?�V'�;�a*9�3�+���θY�q�k{m�{�ʶK���!�����=8�g~�ͻ�^���s�G��x�;���Yא�Mv�j8�x�T��;����'�qMDX��\@x-��r��?KL��k>A��O(�y�d�s�b�[�D�";��T�e��#�,�z�#�sW
�-ӕ�����V�x�8��_7���B4Y _��D9'jI�*��q~Vi9���E�c]nυ�����0*��~�O��b�
�����,���nfJ��}R�89_��X����Yv� ���OOC!�0z����h�I'��Oeu#=((��n���hH�	5�R��L����4�[��	��)�N�r�'��k��Ҁm%B5��w�C�?]���.�'i���-ޢ�[( 1�WG���R�	N_>:�o�w�H���7%���I<�K+������;�na���))�v�D�a<o�<�њZSc���Б7��1%`s�d-������uR=��1(�*2��Mr���36�\t��*]��������O�E"�k���!g|��
�N���l� �mIߨ��N�9H�ة�Ҟ2y��6�հn��'����I��7�����9�>f>�1w$D`^O��!���q�^���~T�B�\��G�]4�\B�`�"]~�
�؝Vf�_"h��(v���m�s�����iL���Y?�9��J�u���x�~�+�1psQp�䣙h=��c�ut��i��ڏqes��mU���SMۨ��ĦX�����!��BuЍ=)3	��� ��`��.Ǝs��.Ӽ�)��\Z�E��W�4�O�wq3Ȣ��&�&3^H��#��R|O�Z=ɣ��ق�%�C����<�,ibd��}�� �YO[~@J�j߰?~��,�8ݯ��4f#�E�c'j�t�������F�꟞i�	V�kWòZ&F��,���[#���k+�r�� i-��Q��-k]g�:�ο6k��yg4�t]�E_0mP�y�IZ���"!&�\�����PJ�!:[��2�`W�_����F���e-��N8�g��98�/�P��AF?sY6n\8^�Y�o��I�~ڒ���u�����vt�E�A�7��G���u~��H���|,F��������P]r����9\f��ZAB�GBծ5�V8Z���d5F(q�-uZ�Qq�"��G�����6���)؏����l	�����Z��fۑ��<�9�J8.�]e�?�%�t���n��?�h@����mH>h��Ԩȏ�x2�}���]y�-�7yV�8��B1R'���c&��j_X{$5�j�]ǥg���-��2���Sg\)�!��
5YgA�7S<B"�Wk��E׸��\)����&�W�:w�|���u�m�Nι���`�����fe�܌$��HIX	�i���$� /ꭨ[$�=Z	�>\g��8L/��tW��{�SM��ܞ4���7���R㧅��JZӖ����7��}����j�|�]�E��L(�a.�ZO�&��W7i�ҋ��g6|��qQ���(H�'�寞��Q��H������/��kHm{�;���e���G79����Cox��[I5���M66�kS�d�+N���qO��� Z����R�"f���#�I��j�҅b�," nM M�ڀt'l���[���f�N�_e�̲\�&�,�'k����0>��M�խ:+Q��I���`$l"�L�,�4�����nԡ��J�8���� h&~w1܉N�r���a���E� ��>Gk<vR���D�e�v�:�����ad���|LB�W��+�/(��՟�p��j���Y���YSvfL�盡wy�e��ޜ7to��o��-r�W�7�|W����F0��V���� ���)z3:6�SG�LNh4��	SD�;j�D�:�*I�	dkl����ko- Em�r��8��8�O�����'%~�����ns�8�y�Y8���꜔��U~ ��O��g��@�-��T��U�}��teȞ5����c��J�6.���"�JB��m�g&�	ɢ��j�bA������c��;[���9�9�FH񱀈��j�L)��� ��\5�@?�<l���L�P;H0	�S�PcQ	Q]�u��9�Ύ�J�#oI$����趱:�G��gf�5��V���f��x����BB_�1�U��}>&��$V8��f7�LH��$.T��,�p#�An���[J��n��"Q�6"&��7�5=��C��,�Kׇ�0t��O�!)eyE\��X���9�G�A	��rȩ�&�0��LY>,�F�o�H�����ЗNeA�����)�^n}᥇�9!��3����?�f�x [z��dV�31���@�hH� ��-T%va�Q@��DC�U)���7:l?qb�8���d}X�uy�m����z]Lw>y�Ĳw���8��V�TC��w�sʮ�+��6�Ĵ1ja�(\�h���-��7m�y��5�i��s5�u���
�T�hBS*2z���Ե��tO��,��]Õ�o��=�8mco�1��hM�/x��4G]1�B5D!�/Ŏ��7����-F4>4�&|9u��5�^Xp�t��3�$|/��g�d�#dY��$�]�=B������@`�8©���gE!��f6/]�8N�|զ��1B���<� ���$�-jQ?D]��ذՊ��� �#Ǹ��G0eBܱ�lnLr�M���r B⠨$�^�֤�r�1?�-'��Iئy�e�O�j<tL��M7A�}c�\��msHS�ݨ��D�Y��{y�S��'>��>xTbuC�з=3��q�I�����f���{�F�%����*	ήS�v�:��?���EHNA�F�`�<�sO 
;��#�AQ���7@8�y�X+��'�]�j��oo�q�����|���	3�g}(�߂��ƭL]��������}����� �9�a\�V���8�lM{������oa��wa`s8�r�n��&�퀉�!�C	�IY���bB�|4�h���v���	�m�3��:��9D�����5��6�~�
|�j��nh�g<����x�Tt�?n��s��������~zk����i*�!�賺�l����>��Gb�΢�:��ʦ�v�g�~A��ƾFu?S|Fi �����f�;�|�b��Oyb&�@���:l��yqK2����w@���'�����	�V�Ι`���!c��m�g߃/x^�@|�%�{ɓ%恪q����'�at������+��ȭ��ܾ�I��eq�c[�UU/�p��7�F��2��8�kE^օ����h�Ow�Ο�� ����#�}��!_$�`|�`�=G�5�Z�q܃�O�hB�b��J)!��}a���#~Hɷq^�#��~�D4_g�3dP�!:�6J�#m�؊��̏��B�
��������
NB�@6� �<��
��y�.4�@@4f�>�?�B�  ؟ԭ�6�*��]��M�tD��NZd��<ݟ��m���P����ey�mn'���
�M�ą�:���a�1�{V�Q���M78ɷ�Z���i�H��C��vcs�=�e��<�u���Ky��{
&8`څ�P��𗃯��ܑ�'��{+��!+;w��&r�}p�9�Z��F��D��7S�������a5��TAR�f4�J��#����ѕ�
��\��Y�-�E��'^�|$�:��N`��g�ZqO��q��%���qG愚ք�a��g�X=��K�܊��"/���wI]54��>�/��B���*�Ŕ���C8��]������׾�Q�����B�W+d���H�7*�尵0�n׏ɥ6l/�x�6��s�Za����<�Ϸ4�nz&�yJ����U�u���ȕ��L�+�3K�����pU�oY:�N�WB��ʚd��=%Oi2s� 4#Y�ሻU���!]�Fx�}ajZ���D�m����Q�_��J1�c3��պP�d�V��f��6�B���F�0L�Os*=չ;�0������s�
ڃ��������/F�x��j)d�![��|-�Ĉ��ޱ�<�M���?� �s{P_�³n�;�/�W�v��N�P!�'�T����y�g��D6�vL�{"��Vh���^��y1�O�,R"K�.�\�`1��CX�O��V8��2yԁ��9�	�xYh�t�Դ�A�}�Q k�J���ha2C���U�v�����*�=`����Wa�Q֯:�7|�?R3�s�#�] G��]QW���j,�s�֏�.'�o�='B_ȅ�����(���<����1z$0���+��:���4�oR2��Is�[&piA�@�$�|r�� q��@:��4x�Q� #�V+����ꟲ65r�h[n�[,�>���҃W���.�G6J6U�Cc `)�1�q.�Ié&���$�x�eH�[]��[�w�Mu�m��#�M[�m����/�6�Bb�iQ��e�Cv&7/�"� ; �}�����!�4Le��>��%$�\��Nt^)jSj@�ma�(l�=�(
QR�H�+n��u���ڷ�5ݸh��t}vsY��n�>�
���(&	Hq!i�D����_���@�:m�"6���������S��o^�����~bB-�c���P3�~'?�M�7�δ�Yy���t��9|Dg��߮�ի�O&З+.��cs[1�VR���<�].㪐�h�!�fS>'���_�C(w�W?w��r{Ѭ���l���"%/ 6���_�̨G1_��|�e������%f���bz�̿xv�@U��8�V/w�qj��Ee[�/����,�n��0�K�6�E�oV�,��4�.�o��]̱��i����f+�������->���3���C(�CJ����p1j5�[�z��j�[���H`�k!�\���1q^�.A�W��Ǯ\��ނ)���D��M��hg��#OC��.uk�$<�4O\��R���|u(�H*�Q���&(�`I���+�����V����#���e��z����F_��w;��Z��C��)���ή�!�\`�|������0%齽��}P�x� ��(̤���zë�S����KI�j�,���|A�$)U�J���iX!)"�Pd�G��>�2��4�ʻ��燉|=�B:��	��p��G�T�uI���}�����;���u�"|C��N96���$�S�mTV�^u�Qkm��ۏx������+s��n��`�R�P�����T�����]br�"=� �;��� Ri��w%a�	t�����:c| e����Ӊ�'��A>��bpe�'����U�N(
M�@"q�|t����?��g�\���a}��Y�Ϙ�����Ѣ,��M�K��m�T�5�5N�B~W�D�>�$�F>�S.�l����ri��%����js_k�J�/_�`<�]r�!D�҆�F�G� �����Nz�T�;3V2K�p���z��:Y��m�P)�f+���<���B�sI0fR	kX.�M�c�3f/�2�m:l
�u; �K䌅�{ �>O³� Q�o�v�	T��Q��	������0��(�`����a?�����d�t�iyԎ��}u�߮s-��k(#���n���Z�t�pY<�%^��?�P�@�8/ٷx�㎁�g�����[l������3��ź˼����:�=�-��ؙ�L+J2� �����g�r�S9��uP,diD�Fqp/Eޔ��^Ltq����S%��L�l�Y٦���S��Qs��ed��c���f�Vu��JԻ�m������w�� ���ӝo���k���������(�pe��y��1Y@��:H�F���P�����Ա ��\�i,^���U��G$֔�����b
�H��f	�����o��	{��J����ɂA��+k�L2�qT��Nn�7��݂�)�h9�r��ݷN\aYh�J�s��	sO)[�y�>���.��z4_v�c�������4󨧆J+WJ3�zIn%.F�A���ŏZR��$��\�(�I
�֕jRZ;r��f_��9)Jq��5\�4��1��q�-;���:~���Xr�������b}g�s��(S��)���<�qS)��ﯬ`O�#���h/a,�Ok�0X#ޮ�E�н'z\�ݖ�:qC���ߵ��4�F���+�!��Kw���{D���v�8�ցGDO�*��L+[�̶������D���'dn���ؼ0��I�<4#g=������#�9}�_N�gqΘ��v��3���gl�����m>��zL�"�l�8�\�`�E��Òa!ה�>ڈp_C8LwS����|}9��P�n��q������M=�AJ]ǭ�%�O%�.[@��[2ܕ
�s�OoZ� 	k���zmX���A?0�(B)��#]� ��vr���3M_ȟ��7U�����e;��� �Xˉgnj^c�Y'��ςG��E�/@�R��Y%aIS\-�C!Mok~cw�E��o�x���SF��J�4l��v��$��c�Szx�x\@�U^�����qQ�+ c�ή-'�S�^5�%ǒ�&c+����@�+��T���4a����-�݄a��'< �"��h[���@8���G1�R��Z�U��3�����M�^�e�	I ���Շ],��y01�eUl�K9@�_մ��*��TN���"@]���A�N��BXi?�(1h��6�����G���2�v���~��F�9߈��h��`@� h-!�gq�d�/Y<�B-�FF��[�~@d�%����U��#B�2p��:R��j�zc�5�,�
\ys��Kv��8ޯ��Y�,�X���V���<��&a�z-�� ����t�k�1�6蘢��8Wi�1�����؀���4"u�P�D�s�(9j�s��4\�ݤ�ε������Ɂ���Nyt�}ĥ���3�=8ȇ�53����/A�Q	��"5�c���������ꪬ��S�tgn��B,t�����<V���QO��N�������q�|�Qg/E���S
��O�0�v��z�mD��V�<$���z�bҧ�>9 d�ڐq�KW��%i�	4m�(��?�`)Z!`����G%���M��˃7��g���2���v�HDœ�Z�R3�}��b�vϙc�%V���G�c�tѨ4 s�XKc(�Y=�/�;�����4��O�u�|V��C�nm����G�N�mh���HV�I��ٸ�ǻ��1�T�YbwW��2���}�/�������$�Sʥc��Z��h�|�Jg?'r��<�� w���,�V�x`� ��	��&*L�Cы�i�YO/v�:E7P1��=������ˣ�G+�,���ؤ�OS��3iQ�����rxq=��~d��yɄKip�T��5`.J=�9�2�J�ʞ��2~������vO�X�.A�ު�K�rk��1�ws:�ݞ�o�	�cz�Z��"�iC7��� W� O7�W[s1�A�����PU�v���Q��y;�6+�1�ċPV�9�l]8���F�Yk�OL�(��y9���2II������i�7M�^~��Ե 3K���y�z���7e�ϳiڍޏQO\J�Cu!K���[E�Yn�B�����D.���c�XtǄ�HPC/ ���vX����Og��-v)�v^	�b�@U0����<�`��_��Q�>�b4�S&�^,.���)o��ͤ�GfmĲ����릘r���	Z�%��v�gu廧��e��A�s(2!w��-�@��'M���f+Q���a/�}Ӗ�K��(a=!ʫoZ2���J��� ��\y^�K�*��2:Y��'�kI(��"�&X���2%[��uث7VFo����q����Ȥ�<��uC��	2�`�����p�#%�L�Z�0�[V�l�yN��CV���ts^��WxaF�A�-'�R��Q�$�|iV�'1⿘�M�S���=2��e�B,���[V 6���,��cܐX���'/Ax�$�^���%���(�����ٴZ�L}��v$3X���z%^_�]5ZR�""�?�a�� Q���5ؕ\���k�B�����d��Q,�Tc_a6��8��@2��� Z�S�$���tf3�c��l���;i��f]=����@�����]�AP.�P��Q]��=�@��1�S�ncD�`�,�ŷ��]&�
< ���>\�F?�n�g��]�݅k

��i5��|����`$F�k3�аu�W��������I��+M��S�����0 ����q�=�t{�<v2Q3�b���hI�Ad�ӷ�ō2%"��������o�� �e�vZ�'c��������~�-J�`���YV��x��:U����R3��E��Mi�تȦ���?��YK����b�*!G��c<x�0ZXk8;�b��-���V����np��a�Kvpγf@|X"�3|��:[��i�za��"���J�~3�β��pJ��eu�h;)ꜨA����Έ���N�3���_��E��UU�0��2���^��b�]jE!)�51ՌzA�.t�����*���������YH�̥�����"�?��3M^ɣ�J��c�R&tV����TDgs��V�t�;�m'4�2�=T/�<��s��lz6p���Sqig�q?������n4Sc
�=G�wvH���!CH\�-�8v)K�<N�}+m-d)ɛ7����,P�&���D
:���v%!b�kg�S;�I��H�ֆr�1�]bt�M,ߺ�lJ�/լcΪ��5�<�Jk�AxP��&�'u��N4$�d�4�q�f�*QK��j�U=��"p�$��zkO���Q�4f�\�?�fh��;�ҝ�%8����@	m~����T��gh��D�����ś��?������Yg)26�m��f�ǅ���X��a�S�������|bc~�ZD+�/曀?EJ%�'C�Ch�q�۝)�_���W�d��Q�Z������3�ժ��]�{�dghNM�[��K�;6��>_��L�4�U��x�n����)}؞��4��.������t�u��(��%�r.�i}����bL8\�\\��r���_� �Omp\S7�L��$��ԦjKt��M�,�c{<'OL�O�7"δ�>7�[�����i����$G\T\�4���d}G����(O"�M3��5����߿�����o�9.��GA�M!�-d&�I,��6W�/�vJ�WU��_��Zd�3~<udL?i�ڔ��\_b;�U��Abr����q����$�5?�U���G�h(�ذ� i���f#���W&9{��;Z��vn��O��.�ƽ�B�H�64��%i�蛌ig�O���m|�QYO�l:���E��M��5�ۓ���qY��jg�����HlC�L,zv{�ǳ!v��w�R��q���I�l��͝����-̲b�jm�Y���H��b<�U!��]��2bͭ���Ή
F"H�[5F �;��`�vC;+�?>N�P�g'��e�[�^�鿖�q�UYg�$�d�M�r0���}\+*�P�!0���"��Z<���ٟk�1HV�|�IH�D����N��q��W�CF$�v��fVN�Th���v�Y GL�\r�0�ߠ�Rp����Y&��5��a3W_�/��Fwv��L](-Kv�FjB�� o������v2q�Rh������}:G�I�������g��au�|3Χ%	g!}���^zA�vN��D�sdEV(�m���]�ƶ:��u$i��R�Z�*��H�O�� ���~bNή��q ���>�?RP�5���g�u��T@��Q�.��d�oW�`z�C���Ӥ���=)�cJ�u\b,�b&���u��A�x_�M�O\�����ꕰ'�07`����%|��T�N��(&\�p㽠c`q�nG���r�CQ���6���B�ד���@���
��:�k�*��絘�����T���|RqECٽD�RT8�����ļ��7Q�E��yI�|�i/#,�%�l���!8 
�@wu��*1v�O��%#�����Y�l�����=K��r,��W)���@��Õ�`�3��R�����d��)�M��BKvt�1�WI@Lt�������t�2C�,b�g]��?R}����2���G�ԝ�~|�?��d�ʜQ���Sk���H �;�Ⱦ��,ѲL�5��Q7���W�ư$���W�z�r^��)ZxU�Q����&��������� ���~��Ib8�qm���qSNH�Z�Oښ�H�`��;�u�߿B�n��ݞ�<�S�����$`��b�v=Rk�I�iH�v�<��g��#T
���O��#6�"@6��b5=э4A��˴2�)�<�=ǘ��Z�;�ں/ՙ�����#m㕅
hr����|L�z�I�r6"tt�ץ��_}E��Csĳ�i�-c��BjH!m��	`��O�gꞙ��|26������5dX����k��ն���=t�.L���� ��0��C�	�\W��Z��os�}��U|J�{��]8�ç�Ik�ܓۇ�7h;�F�J��d��®�MX�۽�a@�Ţ�h��^�S��)|z帡2 ��_���}良�a�d����[V>5L��B,��ײ�,����&T��.�+���2Y<�d8{��5� ��&s�6|�T��h�Eo`�K?r��u�O՟�EC,'�n���?M0n.V������ƷQ�ߓ���
&l����N��.�D�Կ3ȓ��>���v�_���fr��;���1c�Ok�y��D	�uf4.�o�FRӭ?wEL)���ںԏi�Kmp�Y�*x��oқ#f���f�uki��6�XJq
��U�g��l�U�ek�~A�@'��{��TJ;oG;G�lO�"�d�b��X�-`�9���_�7�lߍQz����n"��.�n��A�$�`����a�QR��\L�^��Rm�Ȭ���9(%�W�+up�L���S+��^	��Ф�����,=np�Z�����@1�r��(3Dzg[�Z056�Q���o������XV4����
L٥v���� �ʞ�IJ��#W�N��{�ʊ��t*��8q*}=챽�=6aT�V��I����۳��Zy��+�aol�������cR�P��s��=QA̄еq�J-:��T¹^'�
��y�Cs5�&���c^U��	�� k>�Q�Ў�僜K��9��%N �z�Υv(�7�GfZGWM'�7��w��و������z�,w�2I���в�1��Z��E��X��N�b�������u����r�T��1D��v5mlf��dzW���J���ܓ> ?{��$
Δ�;�ϭ��nC�^�Dkd,�'q��}��z�Q�����U�wZ�~^�|��$��8;'[<��#��t���d�;��|�vwE��K;O�#H�Tx�K�ԽqȖy\�QL�,�������D�h6�^_�P��S!�����{�3c�;�O�)G��K����Gd�: ����[s�-�<���I.��B�sj�b6qޜ�^�P�Z%J@�:�q���\6Qߎ���������� S��Y�de���'v�¨�?���M����Z5/%�J^%z�ǶNAӊ���jk�}�3�Ӽid�Ӕ��k�3�~D�T�k��z�X�U6��]��WfS
�ʇW�/�2�%K�h>d84=�!F?��7�d0����~<�u�,F��T��^�R;�!�P8�+�g�����5�G3�����c�$�^�Pdz������b�D�z�-2�G��0](����;%�	�`.F|�m��<�s_�AD�J�\¶��T|���{��֌���_�Z���}8@��ojPiL�ɀaV����6��H��G�/����)���@p��;���@B��c*������o�ni(��z/O��~yu|���>rc6*2\	ftjw,���!h:�����S��b�)�:n��,�p Bw�;�n����r�*9>���Wsq:g!�1�B(gދ����$#���u��\q�&B�����S��?��� ���	6EgN"����[���1	x������ƣ%��D�1��֮�*�5�#��d��d�-��g��ʚ@�$Qkc�,��IC�7�ɞ�G�8���Qr�yN-߮G��(�1e�*����'Y)Ւ߃� ��!'�ܺ㘩�)De��u�M����x���5�R�\#͈�jK���~���Z�;i��VrN6Q�k����_����T��h���������V�1�d������>�/o�A��B��wS����b{�� ���_S�h�����=`m'͐�,;��V���^��!*`�&�t*ɉ=����,Z'7�Ml�c
�N�V����g�\�L�M�T��W��{�: �GJ:����O� �cq*� �A��$�@���,����F �H4|�����w���P�U����B�S�B��f�8�O��b@��@)ݑ_-���5�gxt�	�h�kW���Iv�2���劕��y>%�d�?���6eK��K���BlTD[�I���Q~Vn��1l�H���tS��}
Ŏ��/dQ�wᦠ(t!�M�>�;W��4���Eg.L,�s��R�RhUУ6g��ȑ��������1�ڴW}���2�\�[38�,{m��(���*웮Wd�A7��{<���)�"t�g��.;�k�U��g�y�0ń�:5�7/�ᶱ��b(�>�lvqY�:y�y�j��r�t1̩�h�����_���i�0� ��g)b�Y�ec�� nb�R�}^ݷ��r�hӆes�B�ւ��9H�i�d������wd�%X	��]g=/oڼov�06mg�x�T��;�f�j�2*��}�׷qR`�e�O�\^�r�(�iIf`��.�'K�|骼��"a��+�W/{��n ٮ5�3�9�?�XG���N�e�X�M����ē���H:�\�dJ�i��?��}�:!S����3boL1!^�:��b(Cb�ą�:���̈�ᚪ��LU���+��|�M��!K_S�������MI\���ZAYx�q��TD6얨�/��
�a��KGc�} ~��zA�R�]��Dm�
�PqiJhb�m�*K�� ��m��\W��Y��/��G/Lz�~�rl���RB�u�M�c4C�o8���1���p4\6y�G|g��J
ְ��Jp�$���lf���UK���O�0�x񮏝��x����B�/\�e�#��!/'�gGLK�޲-���Zc���6��|�;4����_���_������&���B�6����!���*p�����T\����{�ء��8�����0@�x���K>��l�7V[r�$+	������l�u#�/UV`��8]�α),�n�5���JQ�~�����F�a���ߕ�RSR�2��,RnE�/�tu��#M�F��*�cI�7f�0A�b��9%`�r�g�w�����#��@a��������n��Ź�>e�@L<�� 1v#:�r��k�[�����&D�!u�r����J�^��'�oo�l�sH��s��Z�:v0��p٥ Sp�J�K9�uH�Ǫ�y	a)Z��T�^,���{G]�ؑ=1���U�ߏ$q�M����>�$�?��AM��+�q�d�q}@�=8��t����^�`ȥ?X����A����ᢼ�.u-��"Ӊ��/)�RS��v��6��)�t��-�ga�Wβ�i�v�l��,�r欣�3���e�5�3)�\3���UY�<c�d�;r�c�x�l�8ɠ3�ǩ?e�Ν��$��}�(bE*'�9Z^��k�5�8�H�
ӹ��e8Z"�>M3��X���*��>H�C���*���Ӌ����k��K�%�*̑���'��1��ߐ`��&G��,E��r�=������,��qY�]ˆ�ho/���#@��)��.�ơi��-&g�/��c������?��
1X��4��:y�L�3l��WA��|q]g�w�EO���}��G�xw���<�d�eS����#+�%�45����?���̍�����@2�L��eK^����Hf3{���ڽ��N�i/R�웿Q>(|W�u�B*£w���nW���r�N���k����L[�}]�� �B�T�]���Aiʧ�_�3�EC]������.����J�͂R\�Tbq��pM%����H��zoz�#��5������wRRt.c�~z�U�<���?Ex��6,�[_� �]�"���n�>i�h���jj�/~��^vm�)���
d ��I��}6����z�8���Pa���^z �ή���E)�ϕS�s�1 �xY�>���\N��N�0d�-p}�e���]x����@��׭'N���w��Y]�'5eQᮕ��"1�Of��[��g���?"�ZH�-{��^ 8�\�ѐv�I͒K]/�Q�r�..i,>�]�Թ|K��ᒺ!3�`�������fdA�F&T�^� ���)*�=���b߳�F�o}�J�B�D)+�څ�����A���]*=�Cp���ys����ّ^��H�բ^�e���)F�zw�W���fTO��Q���AַK��x��<߰���Q*FOe,�������"R(�L�O�P�m� ��A��ׯ|#��l��.<^'�;��q�nx�>���x�1�G���I���ha勸
�Ɨi��F�T
�����%> �d�!�[�O˱��(���U���y�<H��G%��CTjbFrI4PT�?���R��)�r���J���(p��P�"�F�JEO�lXP�AZ�o�ܤ[���f��, ���k���Ϋ��2��4��/3�`n�a��dP�x��k�00	lTB#�Ф$���ғ'��Y@po*�'Qî0�"'7�t��;t���ޓ� �A%!/GZC��RC� H���'�(
>Bđ���;�	����
� °��hitC����_c<������G��ٺ!J�W��+��5��@zO�nh�fL��E|{�Ȳ֖�K���9���cU����u/sx}��z�hkG,G����{�(���t�B�	u2�ϛ���}d����=�t��{�v����wX���%!˚���Qj�/�GI���A�C�5GXt)nYI:'Jx]=�A����Pe�������cX	E�;�<���O汫H�
��}�Z^�qLf�.UU�@�ҢCa�LR�m٭�h[)�M����-�iэ�y�Kq/�w�x���i��߃�lY��Ȝtg569�&a��ې7Y��hK�M���|�H��$�0�R�(x�PS׫�oI)��F�}r�D��Rq�K�15�0BиMhy�O~�l�Pt�{���!�Gr���رMIm��v(�P�|�I��b��cZ7)���WՏ�5!�S({������}_C5��b��Q��P�:�x��21��B��0�,*�]��~Q�����q �]�ʺ��9�99�\�����z���ZZ���P�M0��
bK�{>}���Y��tV)!�JB%��T�⒓x�G��~g�;���fX�H���4��'w�h4��j/I�����Ao��	-���	��
�v𫽿IW�q��_M��-S�K��ށ�A���B�	=���w7���&u�b�����1��bVӊ
k�����K�]#H�ָ�*�ɜ��.N��^$�]�� moBDT?a�ru�"�x�-��_�t4���e'�#�X0+����<�	f:�%�i���t�Y��ج�y+<	s����똽����R���%�w���K+���T��)g.�s�T����C�� ci�f�2�s���gg������\$l�s&T�rh!��;��&"M?+�4��cj�ID.���3�a���g�b�N����G���j��}�r>M�\=�!y�NP����"��� �z���y^��
c�r&(��S�=�(��hQC�%�}��_5�'2���f�J��˵�*��>�~ѷh�z������5�CK/d�a��1W8/�>I�.�m������ָn��B���v��M�kfv�g/��3�����K��	�L+B'��ڥ�7����//���GVJ5�J�Ѕ��!���f����t�r�}#l�u�h�T2�M��C�KZ�n̑�"�z^aq��^⾶�������K�#���y��`!����q�2 �oݣ�$�8V��耚$AS�h�0�D�����Ĉ-9�Y�&ٌ��!�&�3�F+��ǅ}��B�Ƶ�lko�؂��؀��M?���eᶂ<.�Ϗ�ɺ���q���֜����"A1EwU�S�S�֝�B�7Y�0b�_(��Z�b��P�:N\qFY-��Z��LfQw�ɖ"nkk����:K�A�зCd�)��hy�ȇJ���k�*��L܊����4б�&����z�����)O��E�s���nFKw�a��թ?�ΐȸ��nU�t�e$��S�̈��l����c��w6�}Lƥ�6��j]�RZ_�?1@7�!�,7ԏHo���n���pE�6�s
<��c抈�:E���ꧧW�v���Ű��M�b�[|4.�	�j˘�,������yu<�vj#�7���>׀@@����{��ԕ/Z[�.�A�������C��u��՚�+%W��\>��Z\q��.8W�V���%�؟Rn�����V��k��[��Zɹ��7���
�j�| ���7� �����|��`T-�ѣ�p��a<���c5���@���3�!2*K�X�s�W�+4w���~f)m�J'�RJ*,iᬮV������۬Z�;�61�VZ4�Ɯ���0��#���mߺcC�qm.�I=��jJ4�mˆĉպ�J�y��&p��h��Md�g��F��gqO��`�N��)�}U.�jZ��@�ރh��V��.��^�&��C?�ﰜf*>%]�9�FԳ`�hs� 츌Y���8�W��V���7�B�+؅��~l\l�8���L7��)LO`<��O3b���2nٺ����i���yDJ�@S.��w�o�yW
���5e���:���kj:��{Hs׽�X�`�hM����,��-7F��<�,­M6�@~���Ly��-�e�D���-��m���$+W�0O�:��!djD۪)$l��t-�<�6W/�s6�t���D������7\ѳ��EM��k��Tń��j���(�+-�۴ƯpW�������Vۻ�e2��WK��Ʀ?���;R���==�*�|}h���'�wFS<�.dᶿ�po<�������|��nK@1���(�C^�<��Mm���� ��r�u�x,!�ό�B���ס�_P¢t-g�ug�=���?||�ޒO=���#���!64e�?���뵟:�E2@�z�'��`�D�g�N#x�(��G�^g`�1��?�X��sʼ�d�-�+r��kΫ9�c!rtֳ�5ޮ�w(�/�d���� �B��=K٧*��t���/e��������W����J�K��d���n��5�?iE>�ҟ1�)���/P����΂�Q?u6� �R|�c����J�H�+Uz��P��Wʡ��m��Hd���;��G�7v����5��<�-��ʮ����_
�5�oG��6��F�b�r/�&3�v��zd2�0���.u���6|��[���9 �%US7ѥ�ц:��J�y�v�����)n�R�PdCn�+*7�}�}�m$O��<�!�*��K��K�V1lu1�gMZ��!4��0����4<1N�ua	�S�Ԭ���d&u��'�U���w�c���gs�L�
��|�Kz��X�9d��l���Fx}B}=�1�I��/Zm{K�r���J�E� �O ��ވO��i���o�K�ao����^��e5��a�e����K��BV_i^� s���k�̇fj�Q�U�!!�)!^Q�i|V,������,T�t)���Ϫk��Wyі{���w�9Q l҉ct�/\�u���������p7&�x���;(t6H�k��w�9�WR)�����3�txf�?U
A!�WEp�W�y����}�"��t�)����[�i���-�(VCBأiz�w�c>�y�dE1�Ե����ؚ��	ݶ|z�U�9�'��Lɗ��X��	���������}ǌh�ۍ�Qϧ5+Ɓ��48�i�ÙZ�%&��D$��Uѝ�d�\�V�]�H�4<�=���4��7l(�*|�^��
[7V��/�^�]�l���_����Aֺ��
X�:�2�����u��B�r!�TQ׭�(�N0�g�1t�����u�$O>Xa�T�Gp���W�K��j�y�^� mc~|�>X9Ho���aY�{�y�FL>iz
�X��B��������q�?�G�z�D�H��];�P�o ��C(��0�Q�Ʌ���K�[��XA=��S��]�6Ď"'Qn�3&�zZ8'�4r����@�p3g�5b�ấ�w�1�;O